module Saber_win (
    input logic [13:0] Address,
	 input logic left,
    output logic [23:0] CharacterRGB
);

    // Replace the following data with the 16x16 character's RGB values
    logic [23:0] ROM_Data [12511:0] = '{
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'h7F, 8'h7D, 8'h7F},
{8'h7F, 8'h7F, 8'h78},
{8'h7F, 8'h7E, 8'h79},
{8'h7F, 8'h7D, 8'h7F},
{8'h7F, 8'h7C, 8'h82},
{8'h7E, 8'h7C, 8'h82},
{8'h7C, 8'h7B, 8'h7B},
{8'h96, 8'h95, 8'h8F},
{8'h81, 8'h80, 8'h79},
{8'h80, 8'h7D, 8'h88},
{8'h7F, 8'h7D, 8'h82},
{8'h7C, 8'h7A, 8'h79},
{8'h7E, 8'h7B, 8'h80},
{8'h7C, 8'h78, 8'h84},
{8'h78, 8'h76, 8'h7E},
{8'h7E, 8'h7E, 8'h77},
{8'h82, 8'h83, 8'h70},
{8'h7F, 8'h7D, 8'h86},
{8'h7E, 8'h7D, 8'h82},
{8'h7E, 8'h7F, 8'h79},
{8'h7E, 8'h80, 8'h74},
{8'h7F, 8'h80, 8'h77},
{8'h7E, 8'h7E, 8'h7F},
{8'h7E, 8'h7B, 8'h88},
{8'h7D, 8'h79, 8'h8D},
{8'h79, 8'h80, 8'h7F},
{8'h7C, 8'h83, 8'h81},
{8'h7D, 8'h81, 8'h82},
{8'h7B, 8'h7D, 8'h80},
{8'h7E, 8'h7D, 8'h82},
{8'h7D, 8'h7A, 8'h81},
{8'h81, 8'h7C, 8'h84},
{8'h86, 8'h80, 8'h88},
{8'h7E, 8'h7D, 8'h83},
{8'h7E, 8'h7D, 8'h82},
{8'h7E, 8'h7D, 8'h82},
{8'h7E, 8'h7D, 8'h83},
{8'h80, 8'h7F, 8'h85},
{8'h7E, 8'h7D, 8'h83},
{8'h7E, 8'h7D, 8'h82},
{8'h7F, 8'h7E, 8'h83},
{8'h7C, 8'h7A, 8'h7B},
{8'h80, 8'h7F, 8'h7D},
{8'h81, 8'h84, 8'h7C},
{8'h7A, 8'h7F, 8'h76},
{8'h7B, 8'h7E, 8'h7B},
{8'h7A, 8'h7A, 8'h85},
{8'h81, 8'h7C, 8'h95},
{8'h7E, 8'h76, 8'h98},
{8'h85, 8'h79, 8'h88},
{8'h7F, 8'h7E, 8'h88},
{8'h76, 8'h7F, 8'h87},
{8'h74, 8'h7B, 8'h83},
{8'h7F, 8'h7A, 8'h85},
{8'h84, 8'h7A, 8'h83},
{8'h81, 8'h7C, 8'h81},
{8'h7C, 8'h7F, 8'h7F},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'h7F, 8'h7E, 8'h7A},
{8'h7F, 8'h7E, 8'h7C},
{8'h7F, 8'h7D, 8'h81},
{8'h7F, 8'h7C, 8'h83},
{8'h7E, 8'h7C, 8'h82},
{8'h7B, 8'h79, 8'h7B},
{8'h9B, 8'h9A, 8'h96},
{8'h85, 8'h85, 8'h7E},
{8'h7D, 8'h7B, 8'h7F},
{8'h7A, 8'h79, 8'h74},
{8'h7B, 8'h7C, 8'h6E},
{8'h85, 8'h85, 8'h7A},
{8'h89, 8'h88, 8'h87},
{8'h96, 8'h94, 8'h97},
{8'h87, 8'h86, 8'h82},
{8'h7F, 8'h7F, 8'h73},
{8'h7E, 8'h7D, 8'h81},
{8'h7E, 8'h7E, 8'h81},
{8'h7F, 8'h7E, 8'h7E},
{8'h7F, 8'h7E, 8'h7B},
{8'h7F, 8'h7E, 8'h7C},
{8'h7F, 8'h7C, 8'h80},
{8'h7F, 8'h7A, 8'h83},
{8'h7E, 8'h79, 8'h84},
{8'h7B, 8'h7E, 8'h7B},
{8'h7F, 8'h82, 8'h7D},
{8'h7E, 8'h7F, 8'h7D},
{8'h80, 8'h7E, 8'h7D},
{8'h80, 8'h7D, 8'h7C},
{8'h80, 8'h7B, 8'h7A},
{8'h81, 8'h7A, 8'h79},
{8'h80, 8'h79, 8'h78},
{8'h7A, 8'h77, 8'h75},
{8'h79, 8'h77, 8'h75},
{8'h79, 8'h77, 8'h75},
{8'h7A, 8'h77, 8'h75},
{8'h7C, 8'h7A, 8'h78},
{8'h7D, 8'h7B, 8'h79},
{8'h7F, 8'h7D, 8'h7B},
{8'h80, 8'h7E, 8'h7D},
{8'h7E, 8'h7A, 8'h86},
{8'h7E, 8'h7C, 8'h85},
{8'h81, 8'h7F, 8'h84},
{8'h7D, 8'h7D, 8'h7D},
{8'h7E, 8'h7F, 8'h7C},
{8'h7D, 8'h7C, 8'h7C},
{8'h81, 8'h7F, 8'h81},
{8'h7F, 8'h7B, 8'h7E},
{8'h86, 8'h79, 8'h7D},
{8'h7F, 8'h7D, 8'h7E},
{8'h79, 8'h7F, 8'h7F},
{8'h7A, 8'h7E, 8'h81},
{8'h82, 8'h7C, 8'h83},
{8'h84, 8'h7A, 8'h83},
{8'h80, 8'h7C, 8'h82},
{8'h7A, 8'h80, 8'h82},
{8'h7E, 8'h7D, 8'h80},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'h7F, 8'h7D, 8'h7D},
{8'hFF, 8'hD7, 8'h00},
{8'h7F, 8'h7D, 8'h81},
{8'h7F, 8'h7C, 8'h83},
{8'h80, 8'h7D, 8'h82},
{8'h7A, 8'h78, 8'h79},
{8'hA3, 8'hA2, 8'h9E},
{8'h89, 8'h88, 8'h82},
{8'h7D, 8'h7D, 8'h75},
{8'h93, 8'h95, 8'h7F},
{8'hC9, 8'hCD, 8'hAA},
{8'hE8, 8'hEB, 8'hCB},
{8'hD2, 8'hD4, 8'hC2},
{8'hBE, 8'hBD, 8'hB9},
{8'hB6, 8'hB4, 8'hB4},
{8'h83, 8'h82, 8'h7F},
{8'h7D, 8'h7D, 8'h7B},
{8'h7E, 8'h7E, 8'h80},
{8'h7F, 8'h7C, 8'h83},
{8'h80, 8'h7C, 8'h85},
{8'h80, 8'h7B, 8'h82},
{8'h81, 8'h7A, 8'h7F},
{8'h80, 8'h79, 8'h77},
{8'h7F, 8'h79, 8'h74},
{8'h81, 8'h7E, 8'h79},
{8'h7E, 8'h7A, 8'h73},
{8'h7E, 8'h79, 8'h71},
{8'h7E, 8'h77, 8'h6E},
{8'h85, 8'h7E, 8'h72},
{8'h86, 8'h7E, 8'h70},
{8'h93, 8'h8C, 8'h7C},
{8'hA8, 8'hA1, 8'h90},
{8'hB2, 8'hAE, 8'h9E},
{8'hB2, 8'hAE, 8'h9E},
{8'hB2, 8'hAE, 8'h9E},
{8'hB2, 8'hAE, 8'h9E},
{8'hA3, 8'h9E, 8'h8E},
{8'h8C, 8'h88, 8'h78},
{8'h7C, 8'h78, 8'h67},
{8'h7A, 8'h76, 8'h68},
{8'h7C, 8'h76, 8'h82},
{8'h7F, 8'h78, 8'h87},
{8'h80, 8'h79, 8'h86},
{8'h85, 8'h7F, 8'h87},
{8'h7E, 8'h7A, 8'h79},
{8'h7C, 8'h79, 8'h6D},
{8'h83, 8'h83, 8'h6C},
{8'h83, 8'h81, 8'h67},
{8'h86, 8'h78, 8'h6B},
{8'h79, 8'h74, 8'h67},
{8'h75, 8'h78, 8'h6D},
{8'h81, 8'h82, 8'h7B},
{8'h84, 8'h7B, 8'h7D},
{8'h84, 8'h7A, 8'h81},
{8'h7E, 8'h7D, 8'h85},
{8'h77, 8'h80, 8'h87},
{8'h7E, 8'h7D, 8'h81},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'h7E, 8'h7C, 8'h7F},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'h7E, 8'h7C, 8'h7F},
{8'h7F, 8'h7D, 8'h7F},
{8'h7E, 8'h7C, 8'h7E},
{8'h7E, 8'h7D, 8'h7D},
{8'h7E, 8'h7C, 8'h7C},
{8'h7F, 8'h7E, 8'h7B},
{8'h77, 8'h77, 8'h71},
{8'hA3, 8'hA3, 8'h9B},
{8'h87, 8'h87, 8'h7C},
{8'h9C, 8'h9E, 8'h89},
{8'hF0, 8'hF5, 8'hCF},
{8'hF5, 8'hFC, 8'hC8},
{8'hE6, 8'hEC, 8'hBC},
{8'h8D, 8'h90, 8'h73},
{8'h7C, 8'h7B, 8'h73},
{8'h81, 8'h7F, 8'h82},
{8'h80, 8'h7E, 8'h83},
{8'h7E, 8'h7E, 8'h7A},
{8'h7F, 8'h7D, 8'h7F},
{8'h81, 8'h7D, 8'h87},
{8'h81, 8'h79, 8'h88},
{8'h82, 8'h79, 8'h85},
{8'h82, 8'h79, 8'h79},
{8'h87, 8'h7E, 8'h71},
{8'h8C, 8'h84, 8'h6E},
{8'h95, 8'h8B, 8'h80},
{8'h98, 8'h8D, 8'h81},
{8'h98, 8'h8E, 8'h7E},
{8'hBB, 8'hB4, 8'hA0},
{8'hDB, 8'hD7, 8'hBF},
{8'hF0, 8'hEC, 8'hD0},
{8'hF4, 8'hF0, 8'hD1},
{8'hF9, 8'hF3, 8'hD2},
{8'hFF, 8'hFD, 8'hE1},
{8'hFF, 8'hFE, 8'hE3},
{8'hFF, 8'hFE, 8'hE2},
{8'hFF, 8'hFF, 8'hE3},
{8'hFF, 8'hFD, 8'hE1},
{8'hFA, 8'hF7, 8'hDC},
{8'hE4, 8'hDF, 8'hC3},
{8'hC3, 8'hBD, 8'hA3},
{8'h99, 8'h96, 8'h8D},
{8'h79, 8'h73, 8'h71},
{8'h84, 8'h79, 8'h7D},
{8'h82, 8'h75, 8'h7B},
{8'hA5, 8'h9A, 8'h9A},
{8'hC2, 8'hBB, 8'hB0},
{8'hD2, 8'hD0, 8'hB7},
{8'hE0, 8'hDF, 8'hC0},
{8'hE7, 8'hDD, 8'hC7},
{8'hD0, 8'hCA, 8'hB3},
{8'hA2, 8'hA3, 8'h8D},
{8'h7E, 8'h7B, 8'h6B},
{8'h85, 8'h79, 8'h73},
{8'h86, 8'h7A, 8'h7D},
{8'h7D, 8'h7D, 8'h84},
{8'h76, 8'h80, 8'h88},
{8'h7E, 8'h7D, 8'h81},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'h7E, 8'h7C, 8'h7F},
{8'h7C, 8'h7A, 8'h7D},
{8'h7D, 8'h7B, 8'h7E},
{8'hFF, 8'hD7, 8'h00},
{8'h7F, 8'h7D, 8'h7F},
{8'h78, 8'h77, 8'h74},
{8'h80, 8'h7F, 8'h79},
{8'h80, 8'h80, 8'h76},
{8'h86, 8'h87, 8'h7A},
{8'h7C, 8'h7D, 8'h6C},
{8'h82, 8'h84, 8'h71},
{8'hB8, 8'hBA, 8'hA7},
{8'hAC, 8'hAD, 8'h99},
{8'hBC, 8'hC0, 8'h9C},
{8'hF2, 8'hF8, 8'hC8},
{8'hEF, 8'hF7, 8'hBD},
{8'hF0, 8'hF5, 8'hC4},
{8'h99, 8'h9B, 8'h81},
{8'h7E, 8'h7D, 8'h78},
{8'h7C, 8'h7A, 8'h80},
{8'h7E, 8'h7C, 8'h82},
{8'h81, 8'h81, 8'h7E},
{8'h7C, 8'h7A, 8'h7B},
{8'h81, 8'h7B, 8'h83},
{8'h83, 8'h7A, 8'h85},
{8'h81, 8'h76, 8'h7B},
{8'h7E, 8'h71, 8'h68},
{8'hDD, 8'hD3, 8'hB9},
{8'hF1, 8'hE8, 8'hC5},
{8'hDC, 8'hCD, 8'hB9},
{8'hE6, 8'hD9, 8'hC5},
{8'hFC, 8'hF5, 8'hDD},
{8'hFF, 8'hFF, 8'hE3},
{8'hFE, 8'hF9, 8'hD8},
{8'hF3, 8'hED, 8'hC8},
{8'hEB, 8'hE3, 8'hBA},
{8'hF5, 8'hEF, 8'hC5},
{8'hFF, 8'hFC, 8'hD7},
{8'hFF, 8'hFF, 8'hDC},
{8'hFF, 8'hFC, 8'hD9},
{8'hF7, 8'hF3, 8'hCF},
{8'hEF, 8'hEB, 8'hC7},
{8'hF0, 8'hEB, 8'hC7},
{8'hFF, 8'hFE, 8'hDB},
{8'hFF, 8'hFF, 8'hDC},
{8'hF9, 8'hF8, 8'hD3},
{8'hD3, 8'hD0, 8'hB2},
{8'h9C, 8'h90, 8'h7D},
{8'hA4, 8'h93, 8'h8A},
{8'hB9, 8'hA7, 8'hA2},
{8'hAF, 8'hA1, 8'h9C},
{8'h9C, 8'h93, 8'h8B},
{8'h9D, 8'h98, 8'h8B},
{8'hB2, 8'hA7, 8'h95},
{8'hD3, 8'hCE, 8'hB7},
{8'hFA, 8'hF9, 8'hE1},
{8'hC3, 8'hBC, 8'hA7},
{8'h81, 8'h70, 8'h65},
{8'h8A, 8'h78, 8'h77},
{8'h83, 8'h80, 8'h83},
{8'h7A, 8'h83, 8'h88},
{8'h7E, 8'h7D, 8'h80},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'h81, 8'h7F, 8'h82},
{8'h7E, 8'h7C, 8'h7F},
{8'hFF, 8'hD7, 8'h00},
{8'h7D, 8'h7B, 8'h7D},
{8'hAA, 8'hAB, 8'h9F},
{8'hD1, 8'hD3, 8'hC1},
{8'hD7, 8'hD9, 8'hC1},
{8'hDF, 8'hE2, 8'hC3},
{8'hD0, 8'hD4, 8'hB1},
{8'hE2, 8'hE5, 8'hC1},
{8'hF2, 8'hF6, 8'hD2},
{8'hEF, 8'hF3, 8'hCF},
{8'hED, 8'hF3, 8'hC4},
{8'hEE, 8'hF6, 8'hC1},
{8'hE9, 8'hF1, 8'hBD},
{8'hC5, 8'hC9, 8'hA5},
{8'hAD, 8'hAE, 8'hA1},
{8'h79, 8'h77, 8'h7C},
{8'h7B, 8'h78, 8'h7F},
{8'h80, 8'h7F, 8'h81},
{8'h7F, 8'h7E, 8'h7F},
{8'h82, 8'h7F, 8'h81},
{8'h85, 8'h80, 8'h80},
{8'h84, 8'h7B, 8'h77},
{8'h82, 8'h77, 8'h68},
{8'h92, 8'h84, 8'h6B},
{8'hEF, 8'hE5, 8'hC0},
{8'hE9, 8'hDC, 8'hB2},
{8'hF5, 8'hE9, 8'hCA},
{8'hFF, 8'hFC, 8'hDD},
{8'hF8, 8'hEF, 8'hCF},
{8'hEE, 8'hE6, 8'hC2},
{8'hF5, 8'hEF, 8'hC8},
{8'hFB, 8'hF9, 8'hCF},
{8'hFE, 8'hFC, 8'hD1},
{8'hFD, 8'hFB, 8'hCF},
{8'hFE, 8'hFD, 8'hD6},
{8'hFF, 8'hFE, 8'hD7},
{8'hFC, 8'hF9, 8'hD3},
{8'hEA, 8'hE4, 8'hBE},
{8'hF0, 8'hED, 8'hC7},
{8'hF9, 8'hF6, 8'hD1},
{8'hFF, 8'hFD, 8'hD9},
{8'hFC, 8'hF9, 8'hD3},
{8'hF8, 8'hF9, 8'hC8},
{8'hF0, 8'hEC, 8'hBC},
{8'hEC, 8'hE2, 8'hBA},
{8'hBC, 8'hAB, 8'h8E},
{8'h82, 8'h6C, 8'h5B},
{8'h85, 8'h72, 8'h6C},
{8'h84, 8'h77, 8'h7A},
{8'h83, 8'h7A, 8'h81},
{8'h7F, 8'h76, 8'h6E},
{8'h7A, 8'h77, 8'h67},
{8'h9B, 8'h99, 8'h85},
{8'hEA, 8'hE4, 8'hCF},
{8'hB8, 8'hA4, 8'h96},
{8'h81, 8'h68, 8'h61},
{8'h86, 8'h7D, 8'h78},
{8'h7E, 8'h82, 8'h80},
{8'h7D, 8'h7C, 8'h7F},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'h80, 8'h7E, 8'h81},
{8'h81, 8'h7F, 8'h82},
{8'h81, 8'h7F, 8'h82},
{8'h7A, 8'h78, 8'h7B},
{8'hAC, 8'hAA, 8'hAC},
{8'hD7, 8'hD9, 8'hC2},
{8'hD2, 8'hD5, 8'hB6},
{8'hF6, 8'hFA, 8'hD3},
{8'hF2, 8'hF8, 8'hC9},
{8'hF1, 8'hF9, 8'hC2},
{8'hEE, 8'hF6, 8'hBF},
{8'hEE, 8'hF4, 8'hC0},
{8'hF1, 8'hF8, 8'hC5},
{8'hEC, 8'hF3, 8'hBE},
{8'hEE, 8'hF5, 8'hC2},
{8'hE3, 8'hE8, 8'hC1},
{8'h81, 8'h82, 8'h71},
{8'h81, 8'h7E, 8'h85},
{8'h7C, 8'h78, 8'h89},
{8'h85, 8'h83, 8'h89},
{8'h80, 8'h7F, 8'h7B},
{8'h7E, 8'h7C, 8'h85},
{8'h7E, 8'h7B, 8'h7D},
{8'h81, 8'h7B, 8'h72},
{8'h86, 8'h7F, 8'h67},
{8'hB0, 8'hA7, 8'h84},
{8'h9B, 8'h8D, 8'h64},
{8'hE2, 8'hD2, 8'hA6},
{8'hFC, 8'hF1, 8'hC5},
{8'hF7, 8'hEF, 8'hC8},
{8'hE9, 8'hDD, 8'hB5},
{8'hDD, 8'hD2, 8'hAA},
{8'hF4, 8'hF0, 8'hC7},
{8'hF5, 8'hF3, 8'hC9},
{8'hF9, 8'hF7, 8'hCD},
{8'hF9, 8'hF8, 8'hCF},
{8'hF9, 8'hF8, 8'hCD},
{8'hFF, 8'hFF, 8'hD9},
{8'hFF, 8'hFE, 8'hD9},
{8'hFB, 8'hF8, 8'hD2},
{8'hFC, 8'hFA, 8'hD6},
{8'hFE, 8'hFC, 8'hD7},
{8'hFF, 8'hFF, 8'hDA},
{8'hFD, 8'hFD, 8'hD9},
{8'hF6, 8'hF4, 8'hCF},
{8'hF6, 8'hF4, 8'hCF},
{8'hE9, 8'hE4, 8'hB9},
{8'hF3, 8'hE9, 8'hB8},
{8'hFF, 8'hF6, 8'hC7},
{8'hBB, 8'hA3, 8'h7F},
{8'h84, 8'h71, 8'h5E},
{8'h88, 8'h7B, 8'h7A},
{8'h80, 8'h76, 8'h81},
{8'h82, 8'h7E, 8'h84},
{8'h7D, 8'h7D, 8'h79},
{8'h7D, 8'h7C, 8'h6E},
{8'h92, 8'h84, 8'h72},
{8'hDD, 8'hC5, 8'hB4},
{8'h93, 8'h76, 8'h68},
{8'h83, 8'h73, 8'h68},
{8'h7B, 8'h79, 8'h6F},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'h80, 8'h7E, 8'h81},
{8'h7D, 8'h7B, 8'h7E},
{8'h7E, 8'h7C, 8'h7F},
{8'h7F, 8'h7D, 8'h81},
{8'hA8, 8'hA7, 8'hA8},
{8'h86, 8'h88, 8'h6F},
{8'hBC, 8'hC0, 8'h9D},
{8'hF3, 8'hF9, 8'hCB},
{8'hE8, 8'hF0, 8'hB8},
{8'hF1, 8'hFA, 8'hBC},
{8'hF0, 8'hF8, 8'hB9},
{8'hEE, 8'hF6, 8'hB8},
{8'hEC, 8'hF5, 8'hB8},
{8'hEE, 8'hF5, 8'hBD},
{8'hED, 8'hF3, 8'hC3},
{8'hDA, 8'hDD, 8'hBE},
{8'h89, 8'h88, 8'h84},
{8'h7D, 8'h79, 8'h8A},
{8'h7D, 8'h78, 8'h8D},
{8'h7D, 8'h7B, 8'h7E},
{8'h79, 8'h79, 8'h6D},
{8'h7B, 8'h79, 8'h80},
{8'h7C, 8'h78, 8'h77},
{8'h7F, 8'h79, 8'h66},
{8'hD9, 8'hD3, 8'hAF},
{8'hF1, 8'hE9, 8'hB9},
{8'hC6, 8'hB9, 8'h87},
{8'hFA, 8'hEB, 8'hBB},
{8'hF1, 8'hDF, 8'hB2},
{8'hEF, 8'hE6, 8'hB9},
{8'hF1, 8'hE7, 8'hBC},
{8'hF8, 8'hF1, 8'hC6},
{8'hEF, 8'hE8, 8'hBE},
{8'hF5, 8'hF2, 8'hCA},
{8'hF2, 8'hEF, 8'hC6},
{8'hEC, 8'hEA, 8'hC3},
{8'hFD, 8'hFD, 8'hD9},
{8'hFF, 8'hFF, 8'hD9},
{8'hFE, 8'hFE, 8'hD9},
{8'hFF, 8'hFF, 8'hDC},
{8'hFD, 8'hFD, 8'hD9},
{8'hFC, 8'hFC, 8'hD7},
{8'hF9, 8'hF9, 8'hD3},
{8'hF6, 8'hF5, 8'hD0},
{8'hF2, 8'hF2, 8'hCF},
{8'hF2, 8'hEF, 8'hD6},
{8'hFF, 8'hFB, 8'hDB},
{8'hF2, 8'hE4, 8'hB7},
{8'hFE, 8'hF6, 8'hC1},
{8'hDD, 8'hCD, 8'h9B},
{8'h98, 8'h7E, 8'h5E},
{8'h8B, 8'h75, 8'h6A},
{8'h82, 8'h7A, 8'h7D},
{8'h7E, 8'h7F, 8'h8C},
{8'h79, 8'h7C, 8'h84},
{8'h7E, 8'h7C, 8'h76},
{8'h84, 8'h76, 8'h66},
{8'hA4, 8'h89, 8'h77},
{8'hB0, 8'h8F, 8'h7E},
{8'h85, 8'h6C, 8'h5C},
{8'h86, 8'h80, 8'h70},
{8'h7F, 8'h7D, 8'h7E},
{8'h7F, 8'h7D, 8'h7F},
{8'hFF, 8'hD7, 8'h00},
{8'h7F, 8'h7D, 8'h81},
{8'h7F, 8'h7D, 8'h81},
{8'hFF, 8'hD7, 8'h00},
{8'h7F, 8'h7D, 8'h7F},
{8'h7F, 8'h7D, 8'h7F},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'h80, 8'h7E, 8'h81},
{8'h80, 8'h7E, 8'h81},
{8'hFF, 8'hD7, 8'h00},
{8'h7B, 8'h78, 8'h80},
{8'h9A, 8'h99, 8'h99},
{8'hA8, 8'hA9, 8'h9A},
{8'hB2, 8'hB5, 8'h97},
{8'hD2, 8'hD8, 8'hAC},
{8'hEA, 8'hF0, 8'hBC},
{8'hEF, 8'hF7, 8'hBD},
{8'hED, 8'hF6, 8'hBA},
{8'hEB, 8'hF1, 8'hC3},
{8'hF1, 8'hF7, 8'hCA},
{8'hCF, 8'hD3, 8'hAE},
{8'h7B, 8'h7D, 8'h69},
{8'h7A, 8'h79, 8'h74},
{8'h79, 8'h78, 8'h73},
{8'h78, 8'h79, 8'h64},
{8'hA1, 8'hA7, 8'h80},
{8'hCF, 8'hD7, 8'hAD},
{8'hB6, 8'hB1, 8'h87},
{8'hB5, 8'h9E, 8'h78},
{8'hDF, 8'hC7, 8'hA1},
{8'hD0, 8'hBC, 8'h92},
{8'hE5, 8'hD8, 8'hAB},
{8'hF0, 8'hE5, 8'hB7},
{8'hFC, 8'hF3, 8'hC5},
{8'hED, 8'hEC, 8'hC4},
{8'hF2, 8'hF1, 8'hC9},
{8'hF3, 8'hE9, 8'hC1},
{8'hF4, 8'hE6, 8'hC1},
{8'hEC, 8'hE3, 8'hBE},
{8'hE0, 8'hD1, 8'hAF},
{8'hFA, 8'hF8, 8'hD6},
{8'hFC, 8'hFC, 8'hDC},
{8'hFF, 8'hFE, 8'hD4},
{8'hFC, 8'hFC, 8'hD1},
{8'hF8, 8'hF7, 8'hCD},
{8'hFD, 8'hFC, 8'hD0},
{8'hFE, 8'hFD, 8'hCF},
{8'hF1, 8'hEB, 8'hBD},
{8'hF8, 8'hF3, 8'hC7},
{8'hF1, 8'hED, 8'hBF},
{8'hEB, 8'hFB, 8'hC4},
{8'hFE, 8'hFC, 8'hD7},
{8'hF9, 8'hE5, 8'hD1},
{8'hF4, 8'hF7, 8'hD3},
{8'hF6, 8'hFD, 8'hC8},
{8'hDA, 8'h98, 8'h73},
{8'hB5, 8'h60, 8'h52},
{8'h83, 8'h80, 8'h6A},
{8'h76, 8'h80, 8'h7B},
{8'h78, 8'h7C, 8'h94},
{8'h7F, 8'h7A, 8'h88},
{8'h7B, 8'h83, 8'h78},
{8'h75, 8'h7F, 8'h77},
{8'h99, 8'h6F, 8'h63},
{8'hA1, 8'h64, 8'h4F},
{8'h86, 8'h7B, 8'h6D},
{8'h7C, 8'h7F, 8'h76},
{8'h7E, 8'h7E, 8'h7C},
{8'h7E, 8'h7D, 8'h82},
{8'h7E, 8'h7C, 8'h88},
{8'h7E, 8'h7C, 8'h88},
{8'h7E, 8'h7D, 8'h82},
{8'h7E, 8'h7E, 8'h7B},
{8'h7E, 8'h7F, 8'h77},
{8'h7F, 8'h7D, 8'h7F},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'h80, 8'h7E, 8'h81},
{8'h7D, 8'h7B, 8'h7E},
{8'hFF, 8'hD7, 8'h00},
{8'h7E, 8'h7C, 8'h7F},
{8'h7B, 8'h79, 8'h7C},
{8'h82, 8'h7F, 8'h89},
{8'h79, 8'h76, 8'h7D},
{8'h7A, 8'h79, 8'h79},
{8'h7F, 8'h80, 8'h76},
{8'h7E, 8'h7F, 8'h6A},
{8'hA9, 8'hAD, 8'h8C},
{8'hF1, 8'hF6, 8'hCD},
{8'hEF, 8'hF5, 8'hC6},
{8'hEF, 8'hF6, 8'hC4},
{8'hEE, 8'hF5, 8'hC3},
{8'hE3, 8'hE9, 8'hBE},
{8'hB7, 8'hBA, 8'hA0},
{8'hAA, 8'hAA, 8'h9E},
{8'hB5, 8'hB5, 8'hA9},
{8'hC6, 8'hC9, 8'hAB},
{8'hEC, 8'hF1, 8'hC4},
{8'hF5, 8'hFD, 8'hCC},
{8'hFC, 8'hF7, 8'hCB},
{8'hBC, 8'hA3, 8'h7C},
{8'h8D, 8'h6D, 8'h46},
{8'hD4, 8'hBD, 8'h93},
{8'hF7, 8'hE9, 8'hBB},
{8'hF2, 8'hE3, 8'hB4},
{8'hE0, 8'hCC, 8'h9F},
{8'hE8, 8'hD9, 8'hB3},
{8'hEE, 8'hEC, 8'hC2},
{8'hDC, 8'hD4, 8'hA7},
{8'hF8, 8'hEB, 8'hC2},
{8'hD0, 8'hB8, 8'h90},
{8'hF4, 8'hF1, 8'hC8},
{8'hFE, 8'hFE, 8'hD8},
{8'hFF, 8'hF6, 8'hD4},
{8'hFC, 8'hFA, 8'hD2},
{8'hEA, 8'hE7, 8'hBD},
{8'hF3, 8'hF1, 8'hC6},
{8'hFE, 8'hFD, 8'hD4},
{8'hFF, 8'hFE, 8'hD3},
{8'hE1, 8'hDC, 8'hAF},
{8'hFA, 8'hF6, 8'hCB},
{8'hF5, 8'hEE, 8'hC1},
{8'hF8, 8'hFC, 8'hCA},
{8'hFF, 8'hFE, 8'hDC},
{8'hFC, 8'hF0, 8'hD9},
{8'hEF, 8'hEE, 8'hCC},
{8'hFA, 8'hFF, 8'hCD},
{8'hF8, 8'hD0, 8'hA4},
{8'hBC, 8'h6F, 8'h57},
{8'h87, 8'h71, 8'h57},
{8'h82, 8'h7F, 8'h76},
{8'h7E, 8'h7D, 8'h93},
{8'h81, 8'h7A, 8'h87},
{8'h78, 8'h7F, 8'h76},
{8'h78, 8'h84, 8'h82},
{8'h91, 8'h6C, 8'h65},
{8'h95, 8'h5E, 8'h4D},
{8'h84, 8'h7B, 8'h74},
{8'h7D, 8'h80, 8'h7B},
{8'h7E, 8'h7E, 8'h7D},
{8'h7E, 8'h7D, 8'h83},
{8'h7E, 8'h7C, 8'h87},
{8'h7E, 8'h7C, 8'h87},
{8'h7E, 8'h7D, 8'h83},
{8'h7E, 8'h7E, 8'h7D},
{8'h7E, 8'h7F, 8'h79},
{8'h7F, 8'h7D, 8'h7F},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'h83, 8'h81, 8'h84},
{8'h80, 8'h7E, 8'h81},
{8'h7F, 8'h7D, 8'h7F},
{8'h81, 8'h7F, 8'h81},
{8'h7C, 8'h7A, 8'h7D},
{8'h7F, 8'h7D, 8'h82},
{8'h80, 8'h7D, 8'h86},
{8'h84, 8'h82, 8'h8A},
{8'h7D, 8'h7B, 8'h7C},
{8'h7A, 8'h7A, 8'h6E},
{8'hC5, 8'hC7, 8'hAE},
{8'hF5, 8'hF9, 8'hD6},
{8'hEF, 8'hF7, 8'hC2},
{8'hF4, 8'hFB, 8'hC5},
{8'hD3, 8'hD9, 8'hA9},
{8'hD5, 8'hD9, 8'hB8},
{8'hF5, 8'hF6, 8'hE4},
{8'hEC, 8'hED, 8'hDA},
{8'hF0, 8'hF3, 8'hCE},
{8'hF0, 8'hF7, 8'hC1},
{8'hF1, 8'hF4, 8'hC2},
{8'hDD, 8'hD1, 8'hA5},
{8'hAF, 8'h94, 8'h6E},
{8'h92, 8'h70, 8'h49},
{8'hF3, 8'hDA, 8'hAE},
{8'hF2, 8'hE1, 8'hB2},
{8'hE8, 8'hD5, 8'hA6},
{8'hE0, 8'hC8, 8'h9B},
{8'hF4, 8'hD5, 8'hB2},
{8'hBE, 8'hAE, 8'h7E},
{8'hEF, 8'hE9, 8'hB5},
{8'hCD, 8'hB1, 8'h81},
{8'hEB, 8'hD3, 8'hA3},
{8'hFD, 8'hFF, 8'hCF},
{8'hFB, 8'hFA, 8'hD0},
{8'hFF, 8'hF6, 8'hD4},
{8'hE2, 8'hDC, 8'hB4},
{8'hE2, 8'hDD, 8'hB3},
{8'hFE, 8'hFC, 8'hD3},
{8'hFF, 8'hFC, 8'hD3},
{8'hF2, 8'hEE, 8'hC6},
{8'hD6, 8'hD1, 8'hA8},
{8'hFD, 8'hF8, 8'hCF},
{8'hF9, 8'hF5, 8'hCC},
{8'hFF, 8'hF9, 8'hD2},
{8'hFB, 8'hFF, 8'hDC},
{8'hF8, 8'hF7, 8'hDB},
{8'hEA, 8'hE0, 8'hBE},
{8'hFF, 8'hFF, 8'hCF},
{8'hFF, 8'hF6, 8'hC1},
{8'hD5, 8'h9A, 8'h76},
{8'hA0, 8'h6E, 8'h4D},
{8'h88, 8'h6F, 8'h62},
{8'h83, 8'h7A, 8'h8A},
{8'h86, 8'h7B, 8'h85},
{8'h7D, 8'h7C, 8'h77},
{8'h7A, 8'h84, 8'h87},
{8'h8D, 8'h74, 8'h72},
{8'h86, 8'h5C, 8'h52},
{8'h7C, 8'h77, 8'h7A},
{8'h7E, 8'h80, 8'h80},
{8'h7D, 8'h7D, 8'h7E},
{8'h7D, 8'h7D, 8'h82},
{8'h7E, 8'h7D, 8'h84},
{8'h7E, 8'h7D, 8'h84},
{8'h7E, 8'h7D, 8'h82},
{8'h7E, 8'h7E, 8'h80},
{8'h7E, 8'h7E, 8'h7D},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'h7E, 8'h7C, 8'h7F},
{8'h80, 8'h7E, 8'h81},
{8'h8D, 8'h8B, 8'h8E},
{8'h91, 8'h8F, 8'h92},
{8'h85, 8'h83, 8'h85},
{8'h79, 8'h7A, 8'h6D},
{8'h8C, 8'h8B, 8'h84},
{8'h80, 8'h7D, 8'h81},
{8'h7B, 8'h78, 8'h81},
{8'h7E, 8'h7B, 8'h81},
{8'h7B, 8'h7A, 8'h73},
{8'h81, 8'h83, 8'h6E},
{8'hDF, 8'hE3, 8'hC1},
{8'hEF, 8'hF6, 8'hC0},
{8'hED, 8'hF5, 8'hBC},
{8'hDE, 8'hE5, 8'hB2},
{8'hB9, 8'hBD, 8'h9A},
{8'hD4, 8'hD6, 8'hC0},
{8'hEA, 8'hEB, 8'hD2},
{8'hED, 8'hF3, 8'hC6},
{8'hF1, 8'hF9, 8'hBD},
{8'hE0, 8'hDC, 8'hAB},
{8'hD8, 8'hC7, 8'h9B},
{8'hC6, 8'hAC, 8'h84},
{8'hCA, 8'hA7, 8'h7D},
{8'hFD, 8'hEC, 8'hBE},
{8'hFD, 8'hF2, 8'hC1},
{8'hF9, 8'hE7, 8'hB7},
{8'hF6, 8'hD8, 8'hAC},
{8'hC6, 8'h86, 8'h65},
{8'hD7, 8'hC0, 8'h8E},
{8'hD9, 8'hD0, 8'h96},
{8'hC1, 8'hA2, 8'h6D},
{8'hF9, 8'hE5, 8'hB0},
{8'hF9, 8'hFD, 8'hC4},
{8'hF4, 8'hF4, 8'hC0},
{8'hF1, 8'hD7, 8'hB2},
{8'hC1, 8'hB4, 8'h89},
{8'hFB, 8'hF7, 8'hCD},
{8'hFE, 8'hF9, 8'hD0},
{8'hFD, 8'hF7, 8'hCE},
{8'hCF, 8'hC5, 8'h9C},
{8'hE6, 8'hE1, 8'hBA},
{8'hFD, 8'hFD, 8'hD7},
{8'hFD, 8'hFA, 8'hD2},
{8'hFF, 8'hEE, 8'hD3},
{8'hF2, 8'hFE, 8'hD9},
{8'hF7, 8'hF7, 8'hD7},
{8'hE6, 8'hD2, 8'hB0},
{8'hFD, 8'hFD, 8'hCE},
{8'hFD, 8'hFF, 8'hC6},
{8'hEA, 8'hC4, 8'h93},
{8'hBD, 8'h74, 8'h4A},
{8'h90, 8'h61, 8'h4D},
{8'h85, 8'h75, 8'h7C},
{8'h8A, 8'h7E, 8'h83},
{8'h84, 8'h7D, 8'h7B},
{8'h78, 8'h7F, 8'h89},
{8'h8B, 8'h7E, 8'h7F},
{8'h7C, 8'h60, 8'h58},
{8'h72, 8'h71, 8'h7B},
{8'h7B, 8'h7C, 8'h82},
{8'h85, 8'h84, 8'h86},
{8'h80, 8'h80, 8'h81},
{8'h7E, 8'h7E, 8'h7E},
{8'h7D, 8'h7D, 8'h7C},
{8'h7D, 8'h7D, 8'h7E},
{8'h7D, 8'h7D, 8'h7F},
{8'h7E, 8'h7D, 8'h81},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'h8B, 8'h89, 8'h8C},
{8'hA0, 8'h9E, 8'h9F},
{8'hA7, 8'hAA, 8'h92},
{8'hA4, 8'hA5, 8'h91},
{8'hA4, 8'hA5, 8'h98},
{8'h8C, 8'h8B, 8'h85},
{8'h89, 8'h88, 8'h80},
{8'h94, 8'h95, 8'h85},
{8'h9B, 8'h9E, 8'h82},
{8'hD3, 8'hD7, 8'hB4},
{8'hF2, 8'hF9, 8'hC7},
{8'hE9, 8'hF0, 8'hBC},
{8'hED, 8'hF3, 8'hC3},
{8'hD1, 8'hD5, 8'hB3},
{8'hC8, 8'hCA, 8'hB4},
{8'hF3, 8'hF4, 8'hDC},
{8'hED, 8'hF4, 8'hC7},
{8'hF3, 8'hF8, 8'hBD},
{8'hEF, 8'hE7, 8'hB5},
{8'hA4, 8'h8A, 8'h5D},
{8'hA8, 8'h85, 8'h5B},
{8'hF4, 8'hE3, 8'hB8},
{8'hFC, 8'hEE, 8'hBE},
{8'hFC, 8'hEB, 8'hBA},
{8'hE4, 8'hC8, 8'h98},
{8'hB4, 8'h8A, 8'h5E},
{8'hB1, 8'h6D, 8'h48},
{8'hF6, 8'hDF, 8'hAE},
{8'hB0, 8'h97, 8'h5E},
{8'hD2, 8'hB2, 8'h7A},
{8'hFF, 8'hF5, 8'hBC},
{8'hE7, 8'hE0, 8'hA5},
{8'hE9, 8'hDD, 8'hAA},
{8'hBD, 8'h93, 8'h6C},
{8'hE6, 8'hD7, 8'hA9},
{8'hFF, 8'hFC, 8'hD1},
{8'hEC, 8'hDC, 8'hB2},
{8'hE7, 8'hDA, 8'hB1},
{8'hB0, 8'h9D, 8'h75},
{8'hFA, 8'hF6, 8'hCD},
{8'hFF, 8'hFF, 8'hD6},
{8'hFC, 8'hF8, 8'hD1},
{8'hFD, 8'hE3, 8'hCA},
{8'hF5, 8'hFE, 8'hD8},
{8'hF6, 8'hF7, 8'hD0},
{8'hD3, 8'hB3, 8'h93},
{8'hF7, 8'hF6, 8'hC8},
{8'hF9, 8'hFF, 8'hCB},
{8'hF7, 8'hD6, 8'h9E},
{8'hCE, 8'h7D, 8'h49},
{8'hA1, 8'h60, 8'h45},
{8'h7C, 8'h68, 8'h67},
{8'h82, 8'h78, 8'h76},
{8'h85, 8'h76, 8'h75},
{8'h77, 8'h7B, 8'h87},
{8'h82, 8'h81, 8'h82},
{8'h78, 8'h68, 8'h5F},
{8'h71, 8'h6F, 8'h7A},
{8'h94, 8'h94, 8'h9B},
{8'hE6, 8'hE5, 8'hE6},
{8'hB0, 8'hB2, 8'hAB},
{8'h7B, 8'h7D, 8'h71},
{8'h7F, 8'h81, 8'h76},
{8'h86, 8'h87, 8'h80},
{8'h7C, 8'h7C, 8'h7E},
{8'h7F, 8'h7E, 8'h83},
{8'h80, 8'h7E, 8'h81},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'h80, 8'h7E, 8'h81},
{8'h7C, 8'h7A, 8'h7D},
{8'h7D, 8'h7B, 8'h7F},
{8'h79, 8'h77, 8'h78},
{8'hAA, 8'hAC, 8'h98},
{8'hE8, 8'hEA, 8'hD3},
{8'hAD, 8'hAF, 8'h98},
{8'hC9, 8'hCB, 8'hB3},
{8'hB3, 8'hB6, 8'h9B},
{8'hA7, 8'hAA, 8'h8E},
{8'h9E, 8'hA1, 8'h84},
{8'hA5, 8'hA8, 8'h89},
{8'hE6, 8'hEB, 8'hC2},
{8'hEF, 8'hF5, 8'hC9},
{8'hED, 8'hF2, 8'hCB},
{8'hF1, 8'hF3, 8'hD9},
{8'hF1, 8'hF1, 8'hE3},
{8'hF5, 8'hF6, 8'hE3},
{8'hED, 8'hF3, 8'hCB},
{8'hEC, 8'hF2, 8'hBA},
{8'hFA, 8'hEA, 8'hB8},
{8'h96, 8'h75, 8'h47},
{8'hBF, 8'hA0, 8'h75},
{8'hF5, 8'hDE, 8'hB1},
{8'hE9, 8'hD0, 8'h9F},
{8'hD3, 8'hBB, 8'h88},
{8'hA6, 8'h7F, 8'h4D},
{8'hA0, 8'h6E, 8'h40},
{8'hDF, 8'hAD, 8'h82},
{8'hDC, 8'hB0, 8'h83},
{8'hA6, 8'h73, 8'h41},
{8'hDF, 8'hC0, 8'h88},
{8'hF1, 8'hDD, 8'hA5},
{8'hDD, 8'hBB, 8'h89},
{8'hBE, 8'h97, 8'h6B},
{8'hCA, 8'hAA, 8'h7E},
{8'hFF, 8'hF6, 8'hC4},
{8'hE5, 8'hCC, 8'h9C},
{8'hEB, 8'hD5, 8'hA8},
{8'hC6, 8'hA6, 8'h7C},
{8'hCD, 8'hB8, 8'h8E},
{8'hFF, 8'hFE, 8'hD4},
{8'hFE, 8'hFA, 8'hCF},
{8'hF6, 8'hF3, 8'hC9},
{8'hF1, 8'hDD, 8'hBF},
{8'hFB, 8'hFF, 8'hD5},
{8'hF7, 8'hEF, 8'hC0},
{8'hC2, 8'h9A, 8'h78},
{8'hF6, 8'hF7, 8'hCE},
{8'hF9, 8'hFD, 8'hCF},
{8'hEF, 8'hD3, 8'h99},
{8'hCF, 8'h87, 8'h48},
{8'hAD, 8'h61, 8'h40},
{8'h8C, 8'h7A, 8'h70},
{8'hAA, 8'hA4, 8'h9C},
{8'h99, 8'h86, 8'h82},
{8'h76, 8'h78, 8'h82},
{8'h73, 8'h7A, 8'h74},
{8'h76, 8'h6E, 8'h5E},
{8'h86, 8'h81, 8'h88},
{8'hDB, 8'hDB, 8'hE0},
{8'hFF, 8'hFF, 8'hFC},
{8'hBB, 8'hBE, 8'hAE},
{8'h76, 8'h7A, 8'h62},
{8'hB7, 8'hBB, 8'hA3},
{8'hE3, 8'hE5, 8'hD5},
{8'h9B, 8'h9B, 8'h98},
{8'h7B, 8'h7B, 8'h7F},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'h7D, 8'h7B, 8'h7E},
{8'h80, 8'h7E, 8'h81},
{8'h7E, 8'h7C, 8'h7F},
{8'h75, 8'h73, 8'h76},
{8'hAF, 8'hAE, 8'hAD},
{8'hF9, 8'hF9, 8'hEF},
{8'hD4, 8'hD5, 8'hC0},
{8'h95, 8'h99, 8'h78},
{8'hBA, 8'hBE, 8'h9A},
{8'hA2, 8'hA6, 8'h88},
{8'h7E, 8'h7F, 8'h6A},
{8'hA2, 8'hA3, 8'h93},
{8'hDD, 8'hE1, 8'hC3},
{8'hE7, 8'hEB, 8'hCA},
{8'hE2, 8'hE5, 8'hC9},
{8'hEA, 8'hEB, 8'hDB},
{8'hF7, 8'hF7, 8'hF1},
{8'hF2, 8'hF3, 8'hE7},
{8'hE7, 8'hEB, 8'hCA},
{8'hF2, 8'hF8, 8'hC5},
{8'hE8, 8'hD3, 8'hA2},
{8'h89, 8'h65, 8'h37},
{8'hC7, 8'h9B, 8'h6F},
{8'hCE, 8'hA4, 8'h76},
{8'hB0, 8'h8E, 8'h5C},
{8'hA0, 8'h7E, 8'h4A},
{8'hA9, 8'h7C, 8'h4A},
{8'hC5, 8'h94, 8'h66},
{8'hED, 8'hD8, 8'hA6},
{8'hB4, 8'h70, 8'h48},
{8'hB4, 8'h6A, 8'h41},
{8'hEC, 8'hD3, 8'h9C},
{8'hCD, 8'hB0, 8'h79},
{8'hD9, 8'h96, 8'h6F},
{8'hCE, 8'h8E, 8'h6B},
{8'hEC, 8'hD8, 8'hA8},
{8'hE4, 8'hC8, 8'h90},
{8'hC8, 8'hA3, 8'h6E},
{8'hE6, 8'hC1, 8'h90},
{8'hBF, 8'h92, 8'h64},
{8'hED, 8'hD4, 8'hA8},
{8'hF4, 8'hE8, 8'hBB},
{8'hFC, 8'hF5, 8'hC8},
{8'hE3, 8'hE3, 8'hB4},
{8'hEB, 8'hE7, 8'hC0},
{8'hFF, 8'hFF, 8'hD4},
{8'hF6, 8'hDC, 8'hAB},
{8'hC5, 8'h94, 8'h71},
{8'hF7, 8'hF7, 8'hD4},
{8'hF7, 8'hF6, 8'hD0},
{8'hDE, 8'hC6, 8'h8F},
{8'hCA, 8'h91, 8'h4A},
{8'hB8, 8'h66, 8'h3E},
{8'hCA, 8'hBA, 8'hA9},
{8'hD3, 8'hD1, 8'hC3},
{8'hEE, 8'hE0, 8'hDA},
{8'hB6, 8'hB6, 8'hBD},
{8'hAA, 8'hB7, 8'hAA},
{8'h9D, 8'h99, 8'h7F},
{8'hC6, 8'hBD, 8'hBE},
{8'hFE, 8'hFD, 8'hFE},
{8'hFC, 8'hFD, 8'hF4},
{8'hB6, 8'hB9, 8'hA2},
{8'hAD, 8'hB3, 8'h8F},
{8'hEC, 8'hF2, 8'hCF},
{8'hED, 8'hF0, 8'hD7},
{8'h9A, 8'h9B, 8'h92},
{8'h7D, 8'h7C, 8'h7D},
{8'h80, 8'h7E, 8'h80},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'h7F, 8'h7D, 8'h7F},
{8'h7E, 8'h7C, 8'h7F},
{8'h7F, 8'h7D, 8'h81},
{8'h81, 8'h7F, 8'h82},
{8'h82, 8'h80, 8'h83},
{8'h7D, 8'h7B, 8'h7D},
{8'h7F, 8'h7D, 8'h7C},
{8'h7E, 8'h7D, 8'h7D},
{8'hC6, 8'hC2, 8'hC8},
{8'hFA, 8'hF9, 8'hF5},
{8'hF8, 8'hF8, 8'hE6},
{8'hD7, 8'hDB, 8'hB9},
{8'hDE, 8'hE1, 8'hBE},
{8'hEB, 8'hED, 8'hD3},
{8'hDD, 8'hDD, 8'hD1},
{8'hEE, 8'hEC, 8'hE8},
{8'hEB, 8'hED, 8'hD7},
{8'hE2, 8'hE4, 8'hCC},
{8'hE1, 8'hE2, 8'hCE},
{8'hF0, 8'hF0, 8'hE6},
{8'hFB, 8'hFA, 8'hF8},
{8'hF2, 8'hF1, 8'hEA},
{8'hE7, 8'hEA, 8'hCF},
{8'hED, 8'hF0, 8'hC3},
{8'hD9, 8'hC1, 8'h90},
{8'hA2, 8'h7B, 8'h4D},
{8'hC9, 8'h9F, 8'h73},
{8'hDE, 8'hC2, 8'h93},
{8'hE9, 8'hD6, 8'hA3},
{8'hE7, 8'hCC, 8'h97},
{8'hBB, 8'h8C, 8'h5B},
{8'hED, 8'hCE, 8'h9D},
{8'hD5, 8'hC6, 8'h8E},
{8'h9C, 8'h51, 8'h2A},
{8'hC7, 8'h73, 8'h4F},
{8'hD9, 8'hB9, 8'h86},
{8'hB2, 8'h89, 8'h58},
{8'hE5, 8'h90, 8'h72},
{8'hFC, 8'hB6, 8'h95},
{8'hE1, 8'hD4, 8'h9F},
{8'hB5, 8'h92, 8'h55},
{8'hD8, 8'hA9, 8'h71},
{8'hBC, 8'h8B, 8'h56},
{8'hCA, 8'h9D, 8'h6B},
{8'hF7, 8'hE1, 8'hB3},
{8'hDA, 8'hBF, 8'h8F},
{8'hFE, 8'hFA, 8'hC9},
{8'hCD, 8'hC8, 8'h96},
{8'hE9, 8'hF3, 8'hC2},
{8'hFD, 8'hFD, 8'hC9},
{8'hE7, 8'hC2, 8'h93},
{8'hCD, 8'h97, 8'h74},
{8'hF7, 8'hF6, 8'hD1},
{8'hF4, 8'hEE, 8'hC6},
{8'hD7, 8'hB7, 8'h82},
{8'hCC, 8'h96, 8'h4F},
{8'hAC, 8'h5A, 8'h32},
{8'h96, 8'h86, 8'h74},
{8'hBE, 8'hC0, 8'hB0},
{8'hFF, 8'hF6, 8'hEE},
{8'hF7, 8'hF6, 8'hFA},
{8'hEA, 8'hF8, 8'hEA},
{8'hD4, 8'hD3, 8'hBA},
{8'hF4, 8'hE9, 8'hE7},
{8'hFA, 8'hF9, 8'hFA},
{8'hF9, 8'hFA, 8'hF0},
{8'hD5, 8'hD9, 8'hBC},
{8'hDE, 8'hE6, 8'hBB},
{8'hED, 8'hF5, 8'hC9},
{8'hDA, 8'hDF, 8'hC1},
{8'h82, 8'h85, 8'h77},
{8'h7B, 8'h7B, 8'h7A},
{8'h7E, 8'h7C, 8'h83},
{8'h7F, 8'h7C, 8'h83},
{8'h7F, 8'h7D, 8'h82},
{8'h7F, 8'h7D, 8'h81},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'h7F, 8'h7D, 8'h7F},
{8'h7F, 8'h7D, 8'h7F},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'h80, 8'h7E, 8'h80},
{8'h7E, 8'h7D, 8'h79},
{8'h7F, 8'h7D, 8'h7E},
{8'h7F, 8'h7C, 8'h84},
{8'h7D, 8'h7A, 8'h83},
{8'h84, 8'h82, 8'h85},
{8'h80, 8'h7F, 8'h77},
{8'h7A, 8'h7B, 8'h66},
{8'hB2, 8'hB5, 8'h97},
{8'hF6, 8'hF2, 8'hDC},
{8'hFB, 8'hF9, 8'hE1},
{8'hF4, 8'hF4, 8'hDB},
{8'hED, 8'hEF, 8'hD5},
{8'hF0, 8'hF1, 8'hDC},
{8'hF8, 8'hF6, 8'hE8},
{8'hFB, 8'hF6, 8'hF0},
{8'hF0, 8'hE9, 8'hE6},
{8'hEB, 8'hE9, 8'hD4},
{8'hE1, 8'hDE, 8'hCD},
{8'hE3, 8'hDF, 8'hD6},
{8'hFA, 8'hF5, 8'hF2},
{8'hFE, 8'hFB, 8'hF5},
{8'hF5, 8'hF1, 8'hE2},
{8'hEF, 8'hEE, 8'hD2},
{8'hEB, 8'hEC, 8'hC6},
{8'hBF, 8'hB8, 8'h7F},
{8'h9B, 8'h70, 8'h43},
{8'hEE, 8'hCD, 8'hA7},
{8'hF9, 8'hED, 8'hBD},
{8'hF2, 8'hE3, 8'hB0},
{8'hDC, 8'hBD, 8'h8D},
{8'hC7, 8'hA7, 8'h74},
{8'hFF, 8'hF7, 8'hBC},
{8'hC7, 8'h8E, 8'h5C},
{8'h8C, 8'h47, 8'h17},
{8'hC7, 8'h7D, 8'h53},
{8'hC4, 8'h77, 8'h5A},
{8'hBD, 8'h70, 8'h5E},
{8'hF4, 8'hB7, 8'h9F},
{8'hE1, 8'hAB, 8'h7C},
{8'hB0, 8'h82, 8'h40},
{8'hBF, 8'h8C, 8'h4D},
{8'hE4, 8'h9D, 8'h67},
{8'hEA, 8'hB5, 8'h78},
{8'hCD, 8'hA7, 8'h69},
{8'hDD, 8'hA7, 8'h72},
{8'hDF, 8'hBB, 8'h87},
{8'hF4, 8'hEA, 8'hB3},
{8'hD4, 8'hAE, 8'h7D},
{8'hF4, 8'hF9, 8'hC4},
{8'hF6, 8'hE5, 8'hB9},
{8'hD6, 8'h9E, 8'h7D},
{8'hD5, 8'hA3, 8'h7C},
{8'hF9, 8'hF1, 8'hBA},
{8'hE2, 8'hDD, 8'h9F},
{8'hD0, 8'hA7, 8'h6D},
{8'hE1, 8'h8C, 8'h5E},
{8'hA9, 8'h5D, 8'h41},
{8'h81, 8'h63, 8'h59},
{8'h9F, 8'h9E, 8'h9A},
{8'hFE, 8'hFB, 8'hF1},
{8'hF8, 8'hF1, 8'hEF},
{8'hED, 8'hF0, 8'hFC},
{8'hDF, 8'hDF, 8'hEA},
{8'hF9, 8'hEE, 8'hE9},
{8'hF8, 8'hF3, 8'hFB},
{8'hFA, 8'hFA, 8'hF4},
{8'hEC, 8'hF1, 8'hD2},
{8'hE4, 8'hEE, 8'hBC},
{8'hEA, 8'hF5, 8'hC0},
{8'hC6, 8'hD0, 8'hAA},
{8'h78, 8'h80, 8'h6F},
{8'h77, 8'h7C, 8'h7C},
{8'h78, 8'h76, 8'h87},
{8'h7D, 8'h7A, 8'h8B},
{8'h7E, 8'h7C, 8'h87},
{8'h7B, 8'h7A, 8'h80},
{8'h7E, 8'h7E, 8'h7F},
{8'h7E, 8'h7E, 8'h7E},
{8'h7E, 8'h7E, 8'h7D},
{8'h7E, 8'h7E, 8'h7E},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'h7F, 8'h7D, 8'h7F},
{8'h7E, 8'h7D, 8'h79},
{8'h7E, 8'h7C, 8'h7D},
{8'h7D, 8'h7A, 8'h81},
{8'h7E, 8'h7B, 8'h84},
{8'h78, 8'h76, 8'h79},
{8'h7A, 8'h7A, 8'h72},
{8'h9E, 8'hA0, 8'h8C},
{8'hE7, 8'hE9, 8'hCE},
{8'hF3, 8'hF2, 8'hDF},
{8'hF9, 8'hF7, 8'hE7},
{8'hF6, 8'hF6, 8'hE6},
{8'hF0, 8'hF0, 8'hE2},
{8'hF5, 8'hF5, 8'hEA},
{8'hFC, 8'hFB, 8'hF3},
{8'hFC, 8'hF9, 8'hF3},
{8'hF7, 8'hF3, 8'hEC},
{8'hF3, 8'hF1, 8'hDC},
{8'hE3, 8'hE0, 8'hCF},
{8'hEF, 8'hEB, 8'hE2},
{8'hFE, 8'hFA, 8'hF5},
{8'hFD, 8'hF8, 8'hF2},
{8'hFE, 8'hFC, 8'hED},
{8'hED, 8'hEC, 8'hD3},
{8'hF3, 8'hF3, 8'hD0},
{8'hD8, 8'hCE, 8'h97},
{8'h81, 8'h53, 8'h26},
{8'hAF, 8'h73, 8'h4D},
{8'hC8, 8'hA7, 8'h78},
{8'hC6, 8'hB3, 8'h80},
{8'hCB, 8'hAB, 8'h7C},
{8'hE7, 8'hCF, 8'h9E},
{8'hFF, 8'hF9, 8'hC3},
{8'hAD, 8'h78, 8'h48},
{8'h93, 8'h4F, 8'h23},
{8'hB1, 8'h67, 8'h42},
{8'h82, 8'h3D, 8'h27},
{8'h91, 8'h59, 8'h4C},
{8'h92, 8'h62, 8'h51},
{8'h8B, 8'h53, 8'h34},
{8'h9D, 8'h59, 8'h2E},
{8'hC8, 8'h82, 8'h5A},
{8'hF9, 8'hC0, 8'h93},
{8'hF5, 8'hC0, 8'h92},
{8'hDB, 8'hA4, 8'h75},
{8'hB1, 8'h86, 8'h51},
{8'hF6, 8'hE0, 8'hAC},
{8'hCC, 8'hB0, 8'h7F},
{8'hCF, 8'hBE, 8'h8B},
{8'hF7, 8'hE9, 8'hB6},
{8'hE3, 8'hBD, 8'h90},
{8'hD6, 8'h9E, 8'h75},
{8'hE2, 8'hB4, 8'h86},
{8'hFE, 8'hF3, 8'hBA},
{8'hCE, 8'hB8, 8'h7B},
{8'hC7, 8'h93, 8'h5B},
{8'hD7, 8'h85, 8'h56},
{8'hAB, 8'h62, 8'h41},
{8'h89, 8'h6C, 8'h60},
{8'h6E, 8'h6C, 8'h69},
{8'hDA, 8'hD4, 8'hCB},
{8'hFE, 8'hF3, 8'hF0},
{8'hEB, 8'hED, 8'hF2},
{8'hE5, 8'hE6, 8'hDD},
{8'hFC, 8'hF4, 8'hD5},
{8'hFA, 8'hF6, 8'hF0},
{8'hFA, 8'hF9, 8'hEC},
{8'hEF, 8'hF0, 8'hD6},
{8'hE4, 8'hE8, 8'hC3},
{8'hE7, 8'hEC, 8'hC7},
{8'hB1, 8'hB6, 8'h9B},
{8'h7B, 8'h80, 8'h74},
{8'h8B, 8'h8E, 8'h8B},
{8'h8D, 8'h90, 8'h7E},
{8'h85, 8'h88, 8'h76},
{8'h8A, 8'h8D, 8'h7E},
{8'h82, 8'h84, 8'h79},
{8'h7E, 8'h7F, 8'h79},
{8'h7E, 8'h7E, 8'h7F},
{8'h7E, 8'h7D, 8'h83},
{8'h7E, 8'h7C, 8'h85},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'h7F, 8'h7D, 8'h7F},
{8'h7E, 8'h7D, 8'h7B},
{8'h7C, 8'h7A, 8'h7C},
{8'h9D, 8'h9B, 8'hA1},
{8'hD8, 8'hD5, 8'hDC},
{8'hB5, 8'hB3, 8'hB6},
{8'h93, 8'h92, 8'h8C},
{8'h80, 8'h82, 8'h71},
{8'hCC, 8'hCE, 8'hB8},
{8'hEE, 8'hF0, 8'hE3},
{8'hF7, 8'hF8, 8'hF0},
{8'hF8, 8'hF7, 8'hF3},
{8'hF5, 8'hF3, 8'hF2},
{8'hF9, 8'hF8, 8'hF6},
{8'hFB, 8'hFA, 8'hF5},
{8'hFA, 8'hFA, 8'hF2},
{8'hF8, 8'hF9, 8'hEC},
{8'hEF, 8'hEE, 8'hD9},
{8'hF3, 8'hF0, 8'hDF},
{8'hFD, 8'hF9, 8'hEF},
{8'hFB, 8'hF7, 8'hF0},
{8'hFE, 8'hFA, 8'hF2},
{8'hF6, 8'hF2, 8'hE4},
{8'hE5, 8'hE2, 8'hCD},
{8'hF0, 8'hEE, 8'hD1},
{8'hF7, 8'hED, 8'hB9},
{8'h99, 8'h66, 8'h3E},
{8'h88, 8'h49, 8'h25},
{8'hAF, 8'h8A, 8'h5E},
{8'hE1, 8'hCE, 8'h9D},
{8'hDC, 8'hC1, 8'h94},
{8'hF8, 8'hEA, 8'hBD},
{8'hFE, 8'hFC, 8'hCC},
{8'hBC, 8'h8A, 8'h5D},
{8'h9C, 8'h54, 8'h2F},
{8'h8E, 8'h41, 8'h27},
{8'hBF, 8'h90, 8'h7E},
{8'h91, 8'h86, 8'h78},
{8'h38, 8'h37, 8'h28},
{8'h60, 8'h3F, 8'h2F},
{8'hA2, 8'h5B, 8'h48},
{8'hBF, 8'h71, 8'h5E},
{8'hF4, 8'hCD, 8'hAB},
{8'hE5, 8'hA8, 8'h87},
{8'hCB, 8'h7D, 8'h59},
{8'hC4, 8'hA3, 8'h6E},
{8'hEF, 8'hD6, 8'hA2},
{8'hAB, 8'h7A, 8'h4B},
{8'hEC, 8'hDC, 8'hA6},
{8'hD3, 8'h9B, 8'h6F},
{8'hC1, 8'h83, 8'h55},
{8'hCF, 8'h9D, 8'h6A},
{8'hDE, 8'hB8, 8'h7F},
{8'hFC, 8'hEB, 8'hB1},
{8'hBE, 8'h8A, 8'h54},
{8'hBF, 8'h7C, 8'h4A},
{8'hC1, 8'h75, 8'h45},
{8'hA4, 8'h60, 8'h3A},
{8'h92, 8'h77, 8'h69},
{8'h93, 8'h90, 8'h8F},
{8'hD2, 8'hC7, 8'hC1},
{8'hFE, 8'hEF, 8'hE6},
{8'hED, 8'hED, 8'hE2},
{8'hEB, 8'hEC, 8'hC7},
{8'hF6, 8'hEC, 8'hA8},
{8'hFC, 8'hF8, 8'hDC},
{8'hEF, 8'hEC, 8'hD6},
{8'hF1, 8'hED, 8'hD9},
{8'hF4, 8'hF2, 8'hE0},
{8'hFA, 8'hF8, 8'hE9},
{8'hEE, 8'hEC, 8'hE2},
{8'hE3, 8'hE3, 8'hDD},
{8'hE2, 8'hE1, 8'hDA},
{8'hEA, 8'hF1, 8'hC1},
{8'hE8, 8'hEF, 8'hC1},
{8'hE0, 8'hE6, 8'hC2},
{8'h94, 8'h97, 8'h80},
{8'h7A, 8'h7B, 8'h72},
{8'h7E, 8'h7E, 8'h80},
{8'h7E, 8'h7C, 8'h87},
{8'h7E, 8'h7C, 8'h89},
{8'h7F, 8'h7D, 8'h81},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'h7F, 8'h7D, 8'h7F},
{8'h80, 8'h7E, 8'h7F},
{8'h7D, 8'h7B, 8'h7D},
{8'hA3, 8'hA1, 8'hA6},
{8'hF9, 8'hF6, 8'hFB},
{8'hF5, 8'hF3, 8'hF5},
{8'hEF, 8'hEE, 8'hEA},
{8'hE8, 8'hE7, 8'hDC},
{8'hEF, 8'hEF, 8'hE0},
{8'hEC, 8'hEE, 8'hE7},
{8'hF7, 8'hF8, 8'hF3},
{8'hFC, 8'hF9, 8'hF8},
{8'hFA, 8'hF6, 8'hF5},
{8'hFB, 8'hF6, 8'hF5},
{8'hF9, 8'hF7, 8'hF1},
{8'hF5, 8'hF7, 8'hEC},
{8'hF3, 8'hF6, 8'hE7},
{8'hF4, 8'hF2, 8'hDE},
{8'hFB, 8'hF9, 8'hE9},
{8'hFC, 8'hF9, 8'hED},
{8'hFE, 8'hFC, 8'hF4},
{8'hFF, 8'hFC, 8'hF3},
{8'hFB, 8'hF7, 8'hEB},
{8'hF4, 8'hF2, 8'hE0},
{8'hF2, 8'hF0, 8'hD9},
{8'hDF, 8'hD1, 8'hA5},
{8'hAF, 8'h7C, 8'h59},
{8'h94, 8'h51, 8'h31},
{8'hBF, 8'h99, 8'h6E},
{8'hE6, 8'hD7, 8'hA7},
{8'hE9, 8'hD4, 8'hAA},
{8'hFE, 8'hF6, 8'hCC},
{8'hF7, 8'hF8, 8'hCA},
{8'hC5, 8'h8C, 8'h65},
{8'h9F, 8'h4E, 8'h2F},
{8'h85, 8'h3B, 8'h26},
{8'hDC, 8'hC8, 8'hB7},
{8'h29, 8'h4C, 8'h3B},
{8'h0C, 8'h34, 8'h22},
{8'h16, 8'h20, 8'h11},
{8'h9E, 8'h80, 8'h75},
{8'hDA, 8'hA5, 8'h93},
{8'hCF, 8'hA5, 8'h87},
{8'hCA, 8'h8A, 8'h67},
{8'hE3, 8'h97, 8'h6D},
{8'hE2, 8'hB2, 8'h7D},
{8'hCF, 8'h95, 8'h60},
{8'hB5, 8'h76, 8'h44},
{8'hEE, 8'hC3, 8'h8F},
{8'hD6, 8'h76, 8'h55},
{8'hC9, 8'h80, 8'h55},
{8'hDD, 8'hB3, 8'h79},
{8'hD7, 8'hB3, 8'h76},
{8'hF2, 8'hC2, 8'h8B},
{8'hAE, 8'h5E, 8'h2F},
{8'hB7, 8'h69, 8'h3C},
{8'hB1, 8'h6A, 8'h3C},
{8'h9C, 8'h60, 8'h39},
{8'hDF, 8'hCB, 8'hBC},
{8'hE2, 8'hE3, 8'hE2},
{8'hFD, 8'hF2, 8'hEB},
{8'hF8, 8'hE6, 8'hD9},
{8'hF1, 8'hEF, 8'hD9},
{8'hEA, 8'hED, 8'hB4},
{8'hE1, 8'hD8, 8'h7C},
{8'hEF, 8'hEA, 8'hBF},
{8'hEF, 8'hEA, 8'hCE},
{8'hFB, 8'hF5, 8'hE5},
{8'hFB, 8'hF4, 8'hF0},
{8'hFA, 8'hF3, 8'hF5},
{8'hFD, 8'hF9, 8'hF8},
{8'hFE, 8'hFB, 8'hF5},
{8'hF5, 8'hF3, 8'hE6},
{8'hD5, 8'hDB, 8'hB1},
{8'hC7, 8'hCE, 8'hA6},
{8'hB1, 8'hB5, 8'h99},
{8'h81, 8'h83, 8'h73},
{8'h7D, 8'h7E, 8'h79},
{8'h7E, 8'h7E, 8'h80},
{8'h7E, 8'h7D, 8'h84},
{8'h7E, 8'h7D, 8'h85},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'h7F, 8'h7D, 8'h7F},
{8'h7F, 8'h7D, 8'h7F},
{8'h80, 8'h7E, 8'h80},
{8'h82, 8'h80, 8'h84},
{8'hD1, 8'hCF, 8'hD2},
{8'hF4, 8'hF2, 8'hF3},
{8'hF2, 8'hF1, 8'hEE},
{8'hF7, 8'hF7, 8'hF0},
{8'hF9, 8'hF9, 8'hEF},
{8'hF9, 8'hFB, 8'hF5},
{8'hF4, 8'hF4, 8'hEB},
{8'hF5, 8'hF0, 8'hE3},
{8'hF8, 8'hF1, 8'hE0},
{8'hF2, 8'hEA, 8'hD8},
{8'hF6, 8'hF2, 8'hE1},
{8'hF5, 8'hF5, 8'hE7},
{8'hEC, 8'hEF, 8'hE3},
{8'hEF, 8'hEC, 8'hDB},
{8'hFA, 8'hF8, 8'hE8},
{8'hFB, 8'hF8, 8'hEC},
{8'hFA, 8'hF6, 8'hEC},
{8'hF4, 8'hF0, 8'hE6},
{8'hF0, 8'hEE, 8'hE2},
{8'hF4, 8'hF1, 8'hE4},
{8'hF7, 8'hF4, 8'hE4},
{8'hCF, 8'hC4, 8'hA3},
{8'hC0, 8'h91, 8'h78},
{8'h9F, 8'h5B, 8'h41},
{8'hCA, 8'hA8, 8'h80},
{8'hD6, 8'hC1, 8'h92},
{8'hFB, 8'hE9, 8'hBF},
{8'hFF, 8'hF6, 8'hCC},
{8'hF4, 8'hF6, 8'hC8},
{8'hBF, 8'h7A, 8'h55},
{8'hA4, 8'h50, 8'h32},
{8'hBD, 8'h80, 8'h69},
{8'hCE, 8'hCF, 8'hB9},
{8'h55, 8'h9E, 8'h86},
{8'h38, 8'h8A, 8'h71},
{8'h51, 8'h89, 8'h73},
{8'h9D, 8'hAA, 8'h98},
{8'hFF, 8'hF8, 8'hDB},
{8'hD8, 8'hA8, 8'h89},
{8'hE6, 8'hB6, 8'h89},
{8'hEE, 8'hBB, 8'h84},
{8'hE3, 8'h8F, 8'h5B},
{8'hCE, 8'h77, 8'h41},
{8'hD4, 8'h8D, 8'h55},
{8'hE6, 8'h8D, 8'h60},
{8'hDD, 8'h81, 8'h68},
{8'hE8, 8'hAA, 8'h84},
{8'hFB, 8'hDA, 8'hA5},
{8'hDC, 8'hB5, 8'h7B},
{8'hCE, 8'h84, 8'h55},
{8'hA7, 8'h49, 8'h21},
{8'hAC, 8'h57, 8'h30},
{8'hB2, 8'h70, 8'h45},
{8'hB3, 8'h85, 8'h62},
{8'hD9, 8'hCC, 8'hC0},
{8'hE7, 8'hEA, 8'hEA},
{8'hFD, 8'hF4, 8'hEA},
{8'hFC, 8'hEC, 8'hDB},
{8'hF7, 8'hF4, 8'hDC},
{8'hE9, 8'hEB, 8'hB2},
{8'hE0, 8'hD6, 8'h7B},
{8'hEA, 8'hE5, 8'hBA},
{8'hF9, 8'hF4, 8'hD9},
{8'hFF, 8'hF8, 8'hEB},
{8'hF8, 8'hF1, 8'hF1},
{8'hFB, 8'hF4, 8'hF7},
{8'hFC, 8'hF9, 8'hF5},
{8'hF5, 8'hF3, 8'hE3},
{8'hD5, 8'hD5, 8'hBC},
{8'h9F, 8'hA1, 8'h90},
{8'h7C, 8'h7E, 8'h74},
{8'h78, 8'h79, 8'h75},
{8'h83, 8'h83, 8'h85},
{8'h82, 8'h81, 8'h86},
{8'h80, 8'h80, 8'h83},
{8'h7F, 8'h80, 8'h7F},
{8'h7F, 8'h80, 8'h7C},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'h7E, 8'h7C, 8'h7F},
{8'h7C, 8'h7A, 8'h7D},
{8'hFF, 8'hD7, 8'h00},
{8'h7A, 8'h78, 8'h7B},
{8'h8A, 8'h88, 8'h89},
{8'hD4, 8'hD2, 8'hD2},
{8'hFB, 8'hFA, 8'hF8},
{8'hF4, 8'hF3, 8'hF0},
{8'hF2, 8'hF1, 8'hEE},
{8'hF3, 8'hF2, 8'hEC},
{8'hED, 8'hEA, 8'hD7},
{8'hED, 8'hE5, 8'hC2},
{8'hF4, 8'hE9, 8'hB9},
{8'hF4, 8'hE9, 8'hBA},
{8'hF1, 8'hE9, 8'hC6},
{8'hED, 8'hE9, 8'hD9},
{8'hEA, 8'hE9, 8'hE4},
{8'hE8, 8'hE5, 8'hD6},
{8'hE9, 8'hE5, 8'hD7},
{8'hE7, 8'hE3, 8'hD5},
{8'hEE, 8'hEA, 8'hDE},
{8'hE1, 8'hDD, 8'hD2},
{8'hD9, 8'hD5, 8'hCB},
{8'hE0, 8'hDC, 8'hD3},
{8'hEE, 8'hEA, 8'hE1},
{8'hF0, 8'hEC, 8'hD8},
{8'hB5, 8'h86, 8'h78},
{8'h9E, 8'h5D, 8'h4B},
{8'hD2, 8'hAE, 8'h8A},
{8'hBF, 8'hA8, 8'h79},
{8'hFF, 8'hF0, 8'hC3},
{8'hFF, 8'hF4, 8'hC7},
{8'hF0, 8'hF3, 8'hC1},
{8'hC3, 8'h7A, 8'h52},
{8'hB6, 8'h68, 8'h43},
{8'hE1, 8'hBD, 8'h9B},
{8'hEB, 8'hF6, 8'hDA},
{8'h83, 8'hC4, 8'hAA},
{8'h8E, 8'hE4, 8'hCB},
{8'hA0, 8'hDF, 8'hC3},
{8'hD8, 8'hF3, 8'hD9},
{8'hFC, 8'hFF, 8'hE4},
{8'hF7, 8'hDB, 8'hBC},
{8'hFA, 8'hE1, 8'hB2},
{8'hCC, 8'hA5, 8'h69},
{8'hD9, 8'h84, 8'h51},
{8'hD9, 8'h8C, 8'h59},
{8'hC0, 8'h7E, 8'h48},
{8'hE4, 8'h8D, 8'h67},
{8'h9D, 8'h5F, 8'h4F},
{8'hB8, 8'h8F, 8'h73},
{8'hDD, 8'hC1, 8'h98},
{8'hB4, 8'h7D, 8'h50},
{8'hBF, 8'h6C, 8'h44},
{8'hA2, 8'h42, 8'h20},
{8'hA6, 8'h52, 8'h2F},
{8'hAD, 8'h6C, 8'h47},
{8'h9E, 8'h7D, 8'h65},
{8'h9D, 8'h98, 8'h94},
{8'hBA, 8'hC3, 8'hC3},
{8'hEB, 8'hE4, 8'hD6},
{8'hFD, 8'hEE, 8'hDC},
{8'hF0, 8'hEE, 8'hDC},
{8'hEA, 8'hEC, 8'hC3},
{8'hF3, 8'hE8, 8'hA5},
{8'hF4, 8'hF0, 8'hD2},
{8'hF9, 8'hF6, 8'hE2},
{8'hF8, 8'hF4, 8'hE9},
{8'hF2, 8'hEE, 8'hE8},
{8'hF1, 8'hF0, 8'hE7},
{8'hE7, 8'hE8, 8'hD6},
{8'hE2, 8'hE6, 8'hC6},
{8'hC7, 8'hCD, 8'hA6},
{8'h8C, 8'h8D, 8'h87},
{8'h7B, 8'h7B, 8'h7E},
{8'h7B, 8'h7A, 8'h83},
{8'h7B, 8'h79, 8'h86},
{8'h80, 8'h7E, 8'h89},
{8'h80, 8'h7F, 8'h83},
{8'h7F, 8'h80, 8'h7B},
{8'h7E, 8'h80, 8'h76},
{8'h7F, 8'h7D, 8'h7F},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'h7F, 8'h7D, 8'h82},
{8'h7D, 8'h7B, 8'h7E},
{8'h7D, 8'h7B, 8'h7D},
{8'h7A, 8'h78, 8'h78},
{8'h7E, 8'h7D, 8'h7B},
{8'hBC, 8'hBB, 8'hBA},
{8'hF0, 8'hEF, 8'hF0},
{8'hF3, 8'hF1, 8'hF4},
{8'hEF, 8'hEC, 8'hE1},
{8'hF4, 8'hEE, 8'hCD},
{8'hEE, 8'hE4, 8'hA6},
{8'hE2, 8'hD4, 8'h83},
{8'hE9, 8'hDB, 8'h8C},
{8'hEF, 8'hE3, 8'hAD},
{8'hF5, 8'hED, 8'hDA},
{8'hF8, 8'hF3, 8'hF4},
{8'hE5, 8'hE2, 8'hD5},
{8'hB3, 8'hB0, 8'hA0},
{8'hB1, 8'hAE, 8'h9F},
{8'hA3, 8'hA0, 8'h93},
{8'hE0, 8'hDC, 8'hD1},
{8'hED, 8'hE8, 8'hE0},
{8'hF2, 8'hED, 8'hE7},
{8'hF2, 8'hF0, 8'hEA},
{8'hF7, 8'hF8, 8'hED},
{8'hEB, 8'hC5, 8'hC0},
{8'h91, 8'h53, 8'h46},
{8'h90, 8'h67, 8'h45},
{8'hBC, 8'hA3, 8'h74},
{8'hFF, 8'hF5, 8'hC5},
{8'hFF, 8'hF9, 8'hC9},
{8'hF2, 8'hF1, 8'hBD},
{8'hC2, 8'h7E, 8'h4E},
{8'hB8, 8'h7A, 8'h49},
{8'hEE, 8'hD3, 8'hA4},
{8'hFA, 8'hFA, 8'hDA},
{8'hC2, 8'hDC, 8'hC8},
{8'hA0, 8'hC4, 8'hB2},
{8'h93, 8'hAA, 8'h90},
{8'hEE, 8'hF8, 8'hD9},
{8'hF7, 8'hFA, 8'hE9},
{8'hFA, 8'hF5, 8'hDD},
{8'hF1, 8'hE1, 8'hBC},
{8'hCB, 8'hA2, 8'h73},
{8'hE6, 8'hB6, 8'h83},
{8'hCE, 8'h9C, 8'h6C},
{8'hE6, 8'hB7, 8'h8D},
{8'h96, 8'h6A, 8'h47},
{8'h2F, 8'h23, 8'h16},
{8'h67, 8'h54, 8'h44},
{8'h90, 8'h68, 8'h4D},
{8'h9D, 8'h5B, 8'h3C},
{8'hB7, 8'h60, 8'h40},
{8'h93, 8'h39, 8'h1A},
{8'hAB, 8'h5C, 8'h3C},
{8'h9C, 8'h59, 8'h39},
{8'h7C, 8'h5C, 8'h50},
{8'h63, 8'h68, 8'h69},
{8'h9D, 8'hAE, 8'hAD},
{8'hF4, 8'hF1, 8'hDF},
{8'hFA, 8'hED, 8'hD9},
{8'hED, 8'hEC, 8'hE5},
{8'hEC, 8'hEE, 8'hDE},
{8'hFB, 8'hF0, 8'hCC},
{8'hFA, 8'hF7, 8'hEC},
{8'hF8, 8'hF7, 8'hEF},
{8'hF6, 8'hF6, 8'hEB},
{8'hF2, 8'hF4, 8'hE4},
{8'hE4, 8'hE9, 8'hD0},
{8'hE3, 8'hEA, 8'hC4},
{8'hE5, 8'hF0, 8'hBD},
{8'hEC, 8'hF7, 8'hC1},
{8'hDB, 8'hDE, 8'hC9},
{8'h90, 8'h92, 8'h87},
{8'h7E, 8'h7E, 8'h7D},
{8'h7F, 8'h7E, 8'h87},
{8'h80, 8'h7F, 8'h8A},
{8'h7E, 8'h7D, 8'h83},
{8'h7E, 8'h7E, 8'h7C},
{8'h7D, 8'h7E, 8'h78},
{8'h7F, 8'h7D, 8'h7F},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'h7F, 8'h7D, 8'h82},
{8'h83, 8'h81, 8'h85},
{8'h80, 8'h7E, 8'h7F},
{8'h7D, 8'h7C, 8'h7A},
{8'h7D, 8'h7C, 8'h7B},
{8'h74, 8'h72, 8'h72},
{8'hB2, 8'hB0, 8'hB2},
{8'hF4, 8'hF2, 8'hF4},
{8'hF5, 8'hF0, 8'hE5},
{8'hF3, 8'hEC, 8'hC7},
{8'hEC, 8'hE3, 8'h9C},
{8'hE3, 8'hD7, 8'h7B},
{8'hE0, 8'hD3, 8'h7D},
{8'hF2, 8'hE7, 8'hAE},
{8'hFD, 8'hF5, 8'hE5},
{8'hFE, 8'hF8, 8'hFC},
{8'hFC, 8'hFA, 8'hE9},
{8'hD9, 8'hD7, 8'hC9},
{8'h9F, 8'h9C, 8'h90},
{8'hB1, 8'hB0, 8'h9D},
{8'hF2, 8'hF1, 8'hE0},
{8'hF4, 8'hF0, 8'hEC},
{8'hD6, 8'hD0, 8'hDB},
{8'hA8, 8'hA4, 8'hB4},
{8'h9F, 8'hA4, 8'hB1},
{8'hD6, 8'hB6, 8'hBF},
{8'h6E, 8'h3C, 8'h3B},
{8'h63, 8'h38, 8'h1B},
{8'hCD, 8'hAD, 8'h7E},
{8'hFF, 8'hF5, 8'hCB},
{8'hF9, 8'hEA, 8'hB9},
{8'hF2, 8'hEE, 8'hB1},
{8'hC4, 8'h8E, 8'h57},
{8'hCC, 8'hA2, 8'h68},
{8'hF1, 8'hE3, 8'hAE},
{8'hFB, 8'hF9, 8'hD3},
{8'hF9, 8'hF6, 8'hE3},
{8'hF9, 8'hF1, 8'hE5},
{8'hF7, 8'hF1, 8'hDB},
{8'hFE, 8'hF8, 8'hDA},
{8'hFD, 8'hFA, 8'hF3},
{8'hF7, 8'hFE, 8'hEC},
{8'hFC, 8'hEE, 8'hD3},
{8'hFC, 8'hD9, 8'hB5},
{8'hF1, 8'hE2, 8'hB4},
{8'hF9, 8'hEE, 8'hC3},
{8'hDE, 8'hCC, 8'hAB},
{8'h35, 8'h42, 8'h21},
{8'h00, 8'h13, 8'h07},
{8'h7A, 8'h79, 8'h72},
{8'hDD, 8'hB4, 8'hA3},
{8'hB6, 8'h72, 8'h58},
{8'h9A, 8'h48, 8'h2A},
{8'h9D, 8'h47, 8'h28},
{8'hA7, 8'h58, 8'h3A},
{8'h93, 8'h50, 8'h35},
{8'h7F, 8'h66, 8'h60},
{8'h76, 8'h7C, 8'h7F},
{8'hD7, 8'hE8, 8'hE6},
{8'hF5, 8'hF4, 8'hE2},
{8'hF5, 8'hEA, 8'hD8},
{8'hEE, 8'hEC, 8'hE9},
{8'hEC, 8'hED, 8'hE8},
{8'hEA, 8'hE1, 8'hCE},
{8'hF4, 8'hF3, 8'hEE},
{8'hF7, 8'hF7, 8'hF2},
{8'hF6, 8'hF8, 8'hED},
{8'hF8, 8'hFB, 8'hE8},
{8'hF0, 8'hF7, 8'hD7},
{8'hE2, 8'hED, 8'hBF},
{8'hE4, 8'hF2, 8'hB9},
{8'hDE, 8'hEE, 8'hB0},
{8'hEA, 8'hF2, 8'hC5},
{8'hD3, 8'hD9, 8'hB7},
{8'h81, 8'h84, 8'h71},
{8'h7E, 8'h7F, 8'h7C},
{8'h7E, 8'h7D, 8'h83},
{8'h7E, 8'h7C, 8'h83},
{8'h7D, 8'h7C, 8'h7F},
{8'h7E, 8'h7D, 8'h7D},
{8'h7E, 8'h7D, 8'h81},
{8'h7F, 8'h7D, 8'h82},
{8'h7F, 8'h7D, 8'h82},
{8'h7F, 8'h7D, 8'h82},
{8'h7F, 8'h7D, 8'h81},
{8'hFF, 8'hD7, 8'h00},
{8'h7F, 8'h7D, 8'h7F},
{8'h7F, 8'h7D, 8'h7F},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'h7E, 8'h7C, 8'h81},
{8'h7E, 8'h7C, 8'h80},
{8'h81, 8'h7F, 8'h82},
{8'h7E, 8'h7C, 8'h7E},
{8'h79, 8'h78, 8'h77},
{8'h96, 8'h95, 8'h93},
{8'hEC, 8'hEB, 8'hE8},
{8'hFC, 8'hFB, 8'hF9},
{8'hFA, 8'hF4, 8'hF7},
{8'hF2, 8'hEF, 8'hDD},
{8'hEE, 8'hEF, 8'hC2},
{8'hED, 8'hEF, 8'hBB},
{8'hEB, 8'hEB, 8'hC5},
{8'hEE, 8'hEA, 8'hDB},
{8'hF5, 8'hF0, 8'hF0},
{8'hF7, 8'hF0, 8'hF5},
{8'hF9, 8'hF7, 8'hE5},
{8'hF2, 8'hEF, 8'hEB},
{8'hDF, 8'hDE, 8'hD5},
{8'hAA, 8'hAD, 8'h93},
{8'hA0, 8'hA0, 8'h9D},
{8'h86, 8'h7E, 8'hB4},
{8'h5F, 8'h52, 8'hAC},
{8'h5C, 8'h54, 8'hB2},
{8'h56, 8'h59, 8'hAD},
{8'h7B, 8'h58, 8'h92},
{8'h1F, 8'h10, 8'h49},
{8'h6C, 8'h34, 8'h2A},
{8'hE5, 8'hA7, 8'h6D},
{8'hFC, 8'hFD, 8'hDE},
{8'hE8, 8'hE2, 8'hB1},
{8'hF6, 8'hE7, 8'h9F},
{8'hC1, 8'hA2, 8'h69},
{8'hCF, 8'hC5, 8'h8D},
{8'hE8, 8'hEE, 8'hBD},
{8'hFA, 8'hFA, 8'hD7},
{8'hFF, 8'hF4, 8'hDD},
{8'hFF, 8'hEF, 8'hDD},
{8'hFF, 8'hF5, 8'hDC},
{8'hF9, 8'hFA, 8'hDA},
{8'hFF, 8'hF7, 8'hE8},
{8'hFD, 8'hFB, 8'hE6},
{8'hFA, 8'hFF, 8'hE0},
{8'hFF, 8'hFD, 8'hDB},
{8'hFD, 8'hF9, 8'hD9},
{8'hF3, 8'hF9, 8'hD8},
{8'hAC, 8'hDD, 8'hB3},
{8'h55, 8'hAB, 8'h78},
{8'h27, 8'h6A, 8'h5E},
{8'hA3, 8'hAC, 8'hA7},
{8'hEF, 8'hCB, 8'hBD},
{8'hB6, 8'h87, 8'h60},
{8'h8E, 8'h51, 8'h22},
{8'hAB, 8'h50, 8'h2C},
{8'hA0, 8'h44, 8'h27},
{8'h8E, 8'h53, 8'h34},
{8'h8A, 8'h7E, 8'h6E},
{8'h9F, 8'h9E, 8'h91},
{8'hF7, 8'hF8, 8'hEF},
{8'hF3, 8'hED, 8'hE7},
{8'hF9, 8'hEA, 8'hE4},
{8'hEA, 8'hDB, 8'hCE},
{8'hC5, 8'hBE, 8'hA3},
{8'hB5, 8'hBA, 8'h95},
{8'hCA, 8'hD3, 8'hB5},
{8'hED, 8'hF2, 8'hDD},
{8'hFB, 8'hFB, 8'hEF},
{8'hF5, 8'hF2, 8'hEC},
{8'hF5, 8'hF4, 8'hE9},
{8'hE0, 8'hE3, 8'hCB},
{8'hE1, 8'hE9, 8'hC1},
{8'hE5, 8'hF1, 8'hBD},
{8'hE3, 8'hF3, 8'hB4},
{8'hE9, 8'hF5, 8'hC1},
{8'hA4, 8'hAC, 8'h89},
{8'h75, 8'h78, 8'h69},
{8'h7F, 8'h7D, 8'h7C},
{8'h82, 8'h7D, 8'h83},
{8'h85, 8'h7E, 8'h86},
{8'h81, 8'h79, 8'h82},
{8'h7C, 8'h7B, 8'h85},
{8'h7C, 8'h7C, 8'h87},
{8'h7E, 8'h7D, 8'h88},
{8'h7F, 8'h7D, 8'h88},
{8'h80, 8'h7D, 8'h85},
{8'h80, 8'h7D, 8'h81},
{8'h81, 8'h7C, 8'h7B},
{8'h80, 8'h7C, 8'h79},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'h80, 8'h7E, 8'h81},
{8'h7F, 8'h7D, 8'h82},
{8'h7C, 8'h7A, 8'h7E},
{8'h85, 8'h83, 8'h86},
{8'h7D, 8'h7B, 8'h7D},
{8'h86, 8'h85, 8'h84},
{8'hE0, 8'hDF, 8'hDD},
{8'hFD, 8'hFC, 8'hF9},
{8'hF8, 8'hF7, 8'hF4},
{8'hFA, 8'hF4, 8'hF9},
{8'hF8, 8'hF4, 8'hE9},
{8'hEF, 8'hEF, 8'hCE},
{8'hE9, 8'hE9, 8'hC5},
{8'hFB, 8'hFA, 8'hE1},
{8'hF2, 8'hEE, 8'hE3},
{8'hF5, 8'hF0, 8'hE9},
{8'hFD, 8'hF9, 8'hF3},
{8'hF7, 8'hEF, 8'hF6},
{8'hF2, 8'hEC, 8'hE7},
{8'hD7, 8'hD1, 8'hD4},
{8'h81, 8'h76, 8'h9D},
{8'h5D, 8'h4E, 8'h98},
{8'h5C, 8'h4D, 8'hA1},
{8'h6A, 8'h5C, 8'hAE},
{8'h6A, 8'h5E, 8'hB0},
{8'h7D, 8'h7E, 8'hAD},
{8'h81, 8'h76, 8'hB7},
{8'h51, 8'h3A, 8'h80},
{8'h84, 8'h40, 8'h34},
{8'hD0, 8'hA5, 8'h67},
{8'hF9, 8'hFE, 8'hC4},
{8'hDC, 8'hCF, 8'h89},
{8'hEF, 8'hE5, 8'hBB},
{8'hDB, 8'hAE, 8'h85},
{8'hF3, 8'hDF, 8'hB2},
{8'hEF, 8'hED, 8'hC5},
{8'hFB, 8'hFC, 8'hDD},
{8'hFF, 8'hF8, 8'hE1},
{8'hFF, 8'hF5, 8'hDF},
{8'hFC, 8'hFA, 8'hDC},
{8'hF4, 8'hFF, 8'hDA},
{8'hFA, 8'hFD, 8'hE6},
{8'hF8, 8'hFF, 8'hE3},
{8'hF8, 8'hFF, 8'hDE},
{8'hFF, 8'hFF, 8'hDD},
{8'hF3, 8'hE8, 8'hC9},
{8'hFA, 8'hF8, 8'hDA},
{8'hBB, 8'hD3, 8'hAE},
{8'hA9, 8'hDD, 8'hB5},
{8'h9C, 8'hD2, 8'hBE},
{8'hF3, 8'hF2, 8'hE8},
{8'hF7, 8'hD6, 8'hC6},
{8'h8E, 8'h53, 8'h34},
{8'h97, 8'h52, 8'h2B},
{8'hAD, 8'h54, 8'h31},
{8'hAD, 8'h57, 8'h35},
{8'hA9, 8'h6F, 8'h4B},
{8'h84, 8'h74, 8'h67},
{8'h9D, 8'h98, 8'h8E},
{8'hF5, 8'hF5, 8'hED},
{8'hEE, 8'hE9, 8'hE1},
{8'hF8, 8'hEC, 8'hE2},
{8'hB4, 8'hA5, 8'h91},
{8'hB8, 8'hB2, 8'h8E},
{8'hC3, 8'hCA, 8'h9C},
{8'hC7, 8'hD1, 8'hAE},
{8'hE5, 8'hEA, 8'hD1},
{8'hE6, 8'hE8, 8'hD9},
{8'hF3, 8'hF0, 8'hE9},
{8'hF5, 8'hF2, 8'hE9},
{8'hE1, 8'hE3, 8'hCF},
{8'hA9, 8'hB0, 8'h8D},
{8'hD7, 8'hE3, 8'hB5},
{8'hE5, 8'hF1, 8'hC2},
{8'hEE, 8'hF8, 8'hD1},
{8'hCE, 8'hD3, 8'hBE},
{8'h7D, 8'h7E, 8'h78},
{8'h80, 8'h7E, 8'h83},
{8'h80, 8'h7B, 8'h85},
{8'h81, 8'h7B, 8'h83},
{8'h80, 8'h7A, 8'h81},
{8'h78, 8'h7A, 8'h7B},
{8'h7D, 8'h7F, 8'h7F},
{8'h7F, 8'h80, 8'h82},
{8'h7E, 8'h7E, 8'h80},
{8'h80, 8'h7F, 8'h82},
{8'h80, 8'h7E, 8'h81},
{8'h80, 8'h7D, 8'h80},
{8'h81, 8'h7C, 8'h7F},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'h7F, 8'h7D, 8'h82},
{8'h84, 8'h82, 8'h86},
{8'h82, 8'h80, 8'h83},
{8'h7C, 8'h7A, 8'h7C},
{8'hC2, 8'hC1, 8'hC0},
{8'hFC, 8'hFC, 8'hFA},
{8'hF8, 8'hF7, 8'hF4},
{8'hFB, 8'hFA, 8'hF6},
{8'hFD, 8'hF8, 8'hFC},
{8'hF6, 8'hF2, 8'hED},
{8'hE3, 8'hE1, 8'hD1},
{8'hF6, 8'hF4, 8'hE4},
{8'hF7, 8'hF2, 8'hEA},
{8'hF8, 8'hF3, 8'hED},
{8'hF4, 8'hF0, 8'hE2},
{8'hF0, 8'hEE, 8'hD5},
{8'hFC, 8'hF7, 8'hDA},
{8'hF8, 8'hF3, 8'hE1},
{8'h84, 8'h76, 8'h92},
{8'h3A, 8'h25, 8'h77},
{8'h1C, 8'h0D, 8'h56},
{8'h23, 8'h1A, 8'h3C},
{8'h30, 8'h25, 8'h4C},
{8'h43, 8'h33, 8'h7B},
{8'h63, 8'h58, 8'h83},
{8'h45, 8'h48, 8'h7E},
{8'h52, 8'h37, 8'h58},
{8'h99, 8'h4D, 8'h31},
{8'hBF, 8'h9D, 8'h6F},
{8'hFE, 8'hFF, 8'hCC},
{8'hD8, 8'hCA, 8'h7E},
{8'hEA, 8'hDF, 8'hB6},
{8'hE3, 8'hB1, 8'h91},
{8'hFF, 8'hEB, 8'hCB},
{8'hF1, 8'hEC, 8'hCD},
{8'hFB, 8'hF9, 8'hDF},
{8'hFF, 8'hFC, 8'hE4},
{8'hFF, 8'hFB, 8'hE0},
{8'hFD, 8'hFF, 8'hDD},
{8'hF9, 8'hFF, 8'hDA},
{8'hFB, 8'hFF, 8'hE4},
{8'hFA, 8'hFF, 8'hE1},
{8'hFB, 8'hFF, 8'hDE},
{8'hFE, 8'hFC, 8'hDB},
{8'hF0, 8'hE2, 8'hC5},
{8'hFE, 8'hF7, 8'hDD},
{8'hE7, 8'hE4, 8'hC8},
{8'h99, 8'hA9, 8'h88},
{8'hBE, 8'hDA, 8'hB7},
{8'hFF, 8'hF8, 8'hE1},
{8'hCB, 8'h90, 8'h80},
{8'h90, 8'h43, 8'h2E},
{8'h8F, 8'h40, 8'h24},
{8'hB7, 8'h63, 8'h43},
{8'hC1, 8'h78, 8'h50},
{8'hBF, 8'h92, 8'h66},
{8'h7E, 8'h66, 8'h5D},
{8'h98, 8'h8C, 8'h86},
{8'hE9, 8'hE7, 8'hDF},
{8'hF1, 8'hED, 8'hE3},
{8'hCC, 8'hC0, 8'hB0},
{8'hA8, 8'h9B, 8'h7E},
{8'hBA, 8'hB9, 8'h8B},
{8'hCB, 8'hD5, 8'h9C},
{8'hDE, 8'hE9, 8'hC1},
{8'hF0, 8'hF6, 8'hD9},
{8'hB2, 8'hB4, 8'hA2},
{8'hB5, 8'hB3, 8'hAB},
{8'hE8, 8'hE5, 8'hDD},
{8'hF2, 8'hF3, 8'hE3},
{8'hC6, 8'hCC, 8'hAF},
{8'hBB, 8'hC5, 8'h9F},
{8'hC6, 8'hD1, 8'hAD},
{8'hC8, 8'hD0, 8'hB6},
{8'hB3, 8'hB7, 8'hA9},
{8'h7A, 8'h7C, 8'h79},
{8'h79, 8'h7A, 8'h7C},
{8'h8A, 8'h89, 8'h8B},
{8'h8E, 8'h8C, 8'h8B},
{8'h87, 8'h85, 8'h80},
{8'h80, 8'h87, 8'h77},
{8'h78, 8'h7F, 8'h6F},
{8'h75, 8'h7A, 8'h6D},
{8'h7A, 8'h7C, 8'h73},
{8'h7F, 8'h80, 8'h7D},
{8'h80, 8'h7F, 8'h81},
{8'h80, 8'h7D, 8'h85},
{8'h80, 8'h7C, 8'h85},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'h7E, 8'h7C, 8'h7F},
{8'h7C, 8'h7A, 8'h7F},
{8'h7D, 8'h7B, 8'h7F},
{8'h77, 8'h75, 8'h78},
{8'h9A, 8'h98, 8'h9A},
{8'hF5, 8'hF3, 8'hF3},
{8'hFD, 8'hFD, 8'hFB},
{8'hFA, 8'hFA, 8'hF7},
{8'hF0, 8'hEF, 8'hEB},
{8'hDB, 8'hD6, 8'hD9},
{8'h95, 8'h8F, 8'h8C},
{8'hA5, 8'hA1, 8'h9A},
{8'hFA, 8'hF6, 8'hF4},
{8'hF7, 8'hF0, 8'hF6},
{8'hF6, 8'hF0, 8'hF0},
{8'hF9, 8'hF7, 8'hE7},
{8'hC8, 8'hC7, 8'hA6},
{8'hC2, 8'hBB, 8'h99},
{8'hD8, 8'hD6, 8'hAC},
{8'hCF, 8'hC9, 8'hAD},
{8'h83, 8'h78, 8'h83},
{8'h3B, 8'h30, 8'h51},
{8'h1E, 8'h16, 8'h2E},
{8'h07, 8'h00, 8'h0A},
{8'h25, 8'h1E, 8'h28},
{8'h22, 8'h13, 8'h4B},
{8'h23, 8'h1B, 8'h38},
{8'h41, 8'h20, 8'h10},
{8'h9C, 8'h52, 8'h2A},
{8'hB5, 8'h7F, 8'h66},
{8'hFF, 8'hF6, 8'hD9},
{8'hD9, 8'hC9, 8'h90},
{8'hD6, 8'hC4, 8'h86},
{8'hDC, 8'hB3, 8'h91},
{8'hFC, 8'hE9, 8'hCB},
{8'hF5, 8'hEF, 8'hD3},
{8'hF5, 8'hF3, 8'hD9},
{8'hFF, 8'hFE, 8'hE6},
{8'hFF, 8'hFC, 8'hE1},
{8'hF9, 8'hF1, 8'hD2},
{8'hFA, 8'hEF, 8'hCD},
{8'hF6, 8'hEE, 8'hCF},
{8'hFB, 8'hF4, 8'hD6},
{8'hFF, 8'hFE, 8'hDF},
{8'hFF, 8'hFB, 8'hDC},
{8'hFF, 8'hF8, 8'hDB},
{8'hFB, 8'hF3, 8'hD7},
{8'hFF, 8'hF9, 8'hDC},
{8'hF6, 8'hF7, 8'hD7},
{8'hF3, 8'hF8, 8'hCF},
{8'hF4, 8'hDC, 8'hBC},
{8'h95, 8'h4E, 8'h3D},
{8'h9F, 8'h45, 8'h37},
{8'h89, 8'h32, 8'h1D},
{8'hBA, 8'h6F, 8'h4E},
{8'hC8, 8'h92, 8'h63},
{8'hC5, 8'hA6, 8'h73},
{8'h79, 8'h58, 8'h4F},
{8'h9D, 8'h8B, 8'h85},
{8'hD7, 8'hD3, 8'hC9},
{8'hBD, 8'hBB, 8'hAE},
{8'hB1, 8'hA9, 8'h95},
{8'hB2, 8'hA9, 8'h88},
{8'hAC, 8'hAD, 8'h7C},
{8'hD1, 8'hDB, 8'hA0},
{8'hE8, 8'hF4, 8'hC9},
{8'hBD, 8'hC3, 8'hA4},
{8'h90, 8'h92, 8'h81},
{8'hE6, 8'hE4, 8'hDD},
{8'hAB, 8'hA9, 8'hA3},
{8'hD3, 8'hD4, 8'hC8},
{8'hC4, 8'hCA, 8'hB2},
{8'hC1, 8'hCB, 8'hA9},
{8'hDD, 8'hE5, 8'hC2},
{8'h94, 8'h9B, 8'h7E},
{8'h74, 8'h79, 8'h64},
{8'h79, 8'h7C, 8'h6F},
{8'h7D, 8'h80, 8'h73},
{8'hA0, 8'hA4, 8'h92},
{8'hDD, 8'hE2, 8'hC9},
{8'hD6, 8'hDC, 8'hBE},
{8'hCD, 8'hD8, 8'hB7},
{8'hA3, 8'hAE, 8'h8C},
{8'h91, 8'h9A, 8'h7D},
{8'hA3, 8'hAA, 8'h93},
{8'h8B, 8'h8E, 8'h82},
{8'h80, 8'h81, 8'h80},
{8'h80, 8'h7F, 8'h88},
{8'h80, 8'h7C, 8'h8A},
{8'h7F, 8'h7D, 8'h81},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'h7E, 8'h7C, 8'h81},
{8'h80, 8'h7E, 8'h82},
{8'h7A, 8'h78, 8'h7B},
{8'h91, 8'h8F, 8'h91},
{8'hDE, 8'hDC, 8'hDC},
{8'hC6, 8'hC6, 8'hC3},
{8'h94, 8'h93, 8'h90},
{8'hD3, 8'hD2, 8'hCE},
{8'hD7, 8'hD3, 8'hCF},
{8'h76, 8'h71, 8'h68},
{8'h90, 8'h8C, 8'h83},
{8'hF3, 8'hEE, 8'hEE},
{8'hF8, 8'hF0, 8'hFA},
{8'hF9, 8'hF3, 8'hF8},
{8'hFA, 8'hF8, 8'hEE},
{8'hC1, 8'hC0, 8'hA3},
{8'hAD, 8'hA7, 8'h82},
{8'hAE, 8'hA5, 8'h93},
{8'hDA, 8'hD3, 8'hBF},
{8'hF6, 8'hF4, 8'hD0},
{8'hE3, 8'hDF, 8'hC5},
{8'h8B, 8'h82, 8'h8C},
{8'h1C, 8'h14, 8'h2A},
{8'h26, 8'h20, 8'h30},
{8'h1A, 8'h0D, 8'h49},
{8'h2A, 8'h11, 8'h1D},
{8'h64, 8'h3B, 8'h20},
{8'h84, 8'h41, 8'h2D},
{8'hAD, 8'h5C, 8'h41},
{8'hFC, 8'hE1, 8'hBA},
{8'hE1, 8'hD7, 8'hAF},
{8'hD2, 8'hA4, 8'h69},
{8'hD9, 8'hB8, 8'h8E},
{8'hF4, 8'hE6, 8'hC3},
{8'hFC, 8'hF8, 8'hD8},
{8'hEA, 8'hE9, 8'hCD},
{8'hFD, 8'hFD, 8'hE3},
{8'hFC, 8'hF7, 8'hDD},
{8'hE2, 8'hBE, 8'hA5},
{8'hF4, 8'hBC, 8'hA6},
{8'hEE, 8'hBC, 8'hA2},
{8'hEF, 8'hC3, 8'hA9},
{8'hEA, 8'hCB, 8'hB2},
{8'hF5, 8'hE7, 8'hCA},
{8'hFE, 8'hFE, 8'hDF},
{8'hFB, 8'hFB, 8'hDB},
{8'hF8, 8'hFB, 8'hDA},
{8'hFA, 8'hF9, 8'hD8},
{8'hFF, 8'hFD, 8'hD6},
{8'hC0, 8'hA1, 8'h80},
{8'h8A, 8'h43, 8'h2F},
{8'h9D, 8'h3C, 8'h2D},
{8'h8F, 8'h35, 8'h20},
{8'hBC, 8'h7F, 8'h59},
{8'hD9, 8'hB3, 8'h81},
{8'hCD, 8'hAD, 8'h7A},
{8'h7F, 8'h57, 8'h49},
{8'h93, 8'h7B, 8'h70},
{8'h98, 8'h92, 8'h84},
{8'h8C, 8'h8A, 8'h7B},
{8'hCC, 8'hC5, 8'hB3},
{8'hA7, 8'hA0, 8'h84},
{8'hBC, 8'hBD, 8'h93},
{8'hE7, 8'hF0, 8'hBD},
{8'hDA, 8'hE5, 8'hBC},
{8'h91, 8'h97, 8'h7A},
{8'hC0, 8'hC1, 8'hB2},
{8'hFD, 8'hF9, 8'hF5},
{8'hBA, 8'hB7, 8'hB3},
{8'h81, 8'h82, 8'h76},
{8'hD0, 8'hD4, 8'hBD},
{8'hC9, 8'hD2, 8'hB1},
{8'hB2, 8'hBB, 8'h8E},
{8'hC5, 8'hCD, 8'hA3},
{8'hB3, 8'hBB, 8'h99},
{8'hB8, 8'hC0, 8'hA1},
{8'hD2, 8'hDB, 8'hBA},
{8'hCE, 8'hD9, 8'hB0},
{8'hC4, 8'hD1, 8'h9E},
{8'hE3, 8'hF1, 8'hBA},
{8'hE4, 8'hF2, 8'hC1},
{8'hE3, 8'hF1, 8'hC2},
{8'hE4, 8'hF1, 8'hC5},
{8'hEA, 8'hF4, 8'hD0},
{8'hA8, 8'hAF, 8'h97},
{8'h76, 8'h78, 8'h70},
{8'h7D, 8'h7D, 8'h85},
{8'h7E, 8'h7C, 8'h8B},
{8'h7E, 8'h7C, 8'h81},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'h7F, 8'h7D, 8'h81},
{8'h7D, 8'h7B, 8'h80},
{8'h7D, 8'h7B, 8'h7F},
{8'hFF, 8'hD7, 8'h00},
{8'h7B, 8'h79, 8'h7B},
{8'h7F, 8'h7E, 8'h7D},
{8'h75, 8'h74, 8'h72},
{8'h8F, 8'h8E, 8'h8B},
{8'hEE, 8'hED, 8'hE8},
{8'hEC, 8'hE9, 8'hDB},
{8'hB2, 8'hAF, 8'h9B},
{8'hBE, 8'hBC, 8'hA6},
{8'hF3, 8'hF1, 8'hE5},
{8'hFB, 8'hF6, 8'hFA},
{8'hFF, 8'hFA, 8'hFF},
{8'hFF, 8'hFA, 8'hFE},
{8'hC7, 8'hC3, 8'hBA},
{8'hC3, 8'hBB, 8'hAC},
{8'hE6, 8'hDC, 8'hE6},
{8'hFB, 8'hF4, 8'hF8},
{8'hD5, 8'hD4, 8'hB6},
{8'hCB, 8'hCB, 8'hA9},
{8'h3D, 8'h37, 8'h45},
{8'h19, 8'h0D, 8'h41},
{8'h2D, 8'h22, 8'h5B},
{8'h09, 8'h05, 8'h38},
{8'h19, 8'h0C, 8'h11},
{8'h6A, 8'h43, 8'h2E},
{8'h66, 8'h2E, 8'h2F},
{8'hA4, 8'h53, 8'h2E},
{8'hE3, 8'hBA, 8'h71},
{8'hF5, 8'hF0, 8'hC8},
{8'hC9, 8'h88, 8'h62},
{8'hCB, 8'hA1, 8'h73},
{8'hDA, 8'hBE, 8'h96},
{8'hFF, 8'hF9, 8'hD7},
{8'hEB, 8'hE5, 8'hC6},
{8'hF9, 8'hFA, 8'hDC},
{8'hFB, 8'hF7, 8'hDB},
{8'hED, 8'hC1, 8'hAB},
{8'hFF, 8'hBE, 8'hAD},
{8'hFE, 8'hBE, 8'hA2},
{8'hFE, 8'hC1, 8'hA8},
{8'hE5, 8'hAF, 8'h97},
{8'hE7, 8'hCF, 8'hB2},
{8'hFE, 8'hFF, 8'hE2},
{8'hF6, 8'hFF, 8'hDF},
{8'hF9, 8'hFE, 8'hDB},
{8'hFF, 8'hFF, 8'hDE},
{8'hEC, 8'hE1, 8'hC7},
{8'h90, 8'h75, 8'h5A},
{8'h92, 8'h53, 8'h3C},
{8'h96, 8'h35, 8'h20},
{8'h96, 8'h3F, 8'h21},
{8'hC0, 8'h93, 8'h64},
{8'hEB, 8'hDA, 8'hA5},
{8'hBE, 8'hA2, 8'h73},
{8'h8F, 8'h60, 8'h49},
{8'h9E, 8'h82, 8'h6C},
{8'h8E, 8'h86, 8'h72},
{8'hAD, 8'hAB, 8'h9C},
{8'hBC, 8'hB6, 8'hAA},
{8'hAF, 8'hA8, 8'h98},
{8'hA5, 8'hA4, 8'h8D},
{8'hCC, 8'hD3, 8'hB4},
{8'h9B, 8'hA5, 8'h83},
{8'hD6, 8'hDB, 8'hC3},
{8'hF0, 8'hF1, 8'hE5},
{8'hF8, 8'hF5, 8'hF2},
{8'hE3, 8'hE0, 8'hDC},
{8'h7C, 8'h7D, 8'h70},
{8'h81, 8'h86, 8'h6B},
{8'hBF, 8'hC9, 8'hA4},
{8'hD4, 8'hDD, 8'hAA},
{8'hE3, 8'hEC, 8'hBC},
{8'hE8, 8'hF1, 8'hC7},
{8'hE8, 8'hF3, 8'hCB},
{8'hE6, 8'hF3, 8'hC7},
{8'hE6, 8'hF6, 8'hC1},
{8'hDE, 8'hF1, 8'hB3},
{8'hDE, 8'hF2, 8'hAE},
{8'hDF, 8'hF0, 8'hB7},
{8'hE0, 8'hF1, 8'hBA},
{8'hE3, 8'hF2, 8'hBC},
{8'hE5, 8'hF2, 8'hC2},
{8'h9D, 8'hA7, 8'h84},
{8'h78, 8'h7D, 8'h6D},
{8'h78, 8'h79, 8'h7B},
{8'h7B, 8'h7B, 8'h86},
{8'h7F, 8'h7D, 8'h81},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'h7D, 8'h7B, 8'h80},
{8'h7E, 8'h7C, 8'h80},
{8'h7E, 8'h7C, 8'h7F},
{8'h81, 8'h7F, 8'h81},
{8'h83, 8'h81, 8'h81},
{8'h79, 8'h77, 8'h76},
{8'h9B, 8'h9A, 8'h98},
{8'hED, 8'hEC, 8'hE7},
{8'hEC, 8'hEA, 8'hD4},
{8'hE6, 8'hE6, 8'hC5},
{8'hF4, 8'hF5, 8'hD0},
{8'hF5, 8'hF3, 8'hDA},
{8'hFD, 8'hFA, 8'hF5},
{8'hDA, 8'hD3, 8'hDE},
{8'hA6, 8'h9F, 8'hAC},
{8'hA8, 8'hA0, 8'hAF},
{8'hF1, 8'hE8, 8'hF8},
{8'hFB, 8'hF8, 8'hF1},
{8'hF9, 8'hF8, 8'hDF},
{8'hCE, 8'hCC, 8'hBA},
{8'h9D, 8'h98, 8'hA3},
{8'h5E, 8'h57, 8'h7D},
{8'h80, 8'h78, 8'hA2},
{8'h8C, 8'h83, 8'hB0},
{8'h57, 8'h61, 8'h97},
{8'h2D, 8'h4F, 8'h59},
{8'h86, 8'h70, 8'h41},
{8'hBC, 8'h8E, 8'h7C},
{8'h8E, 8'h54, 8'h3F},
{8'hB1, 8'h88, 8'h40},
{8'hF9, 8'hF4, 8'hBB},
{8'hCD, 8'h99, 8'h6D},
{8'hD6, 8'h94, 8'h65},
{8'hBF, 8'h80, 8'h57},
{8'hFB, 8'hDA, 8'hB8},
{8'hF1, 8'hE6, 8'hC5},
{8'hF6, 8'hF9, 8'hD9},
{8'hFF, 8'hFE, 8'hDF},
{8'hF4, 8'hD1, 8'hB8},
{8'hFB, 8'hB9, 8'hA7},
{8'hFE, 8'hC0, 8'h9C},
{8'hFC, 8'hBC, 8'h9E},
{8'hEF, 8'hBB, 8'hA1},
{8'hFC, 8'hEE, 8'hD0},
{8'hF9, 8'hFF, 8'hDF},
{8'hF7, 8'hFF, 8'hE1},
{8'hFF, 8'hFF, 8'hDE},
{8'hF5, 8'hE1, 8'hC6},
{8'h9E, 8'h8A, 8'h83},
{8'h7E, 8'h6B, 8'h5A},
{8'h72, 8'h3F, 8'h24},
{8'h99, 8'h3C, 8'h20},
{8'hA9, 8'h58, 8'h30},
{8'hD5, 8'hB7, 8'h7F},
{8'hFE, 8'hFC, 8'hC6},
{8'hA0, 8'h82, 8'h57},
{8'h91, 8'h62, 8'h3F},
{8'hD2, 8'hB9, 8'h99},
{8'hCC, 8'hC2, 8'hAB},
{8'hF5, 8'hF5, 8'hE8},
{8'hEC, 8'hE8, 8'hE3},
{8'hEB, 8'hE5, 8'hE3},
{8'hB2, 8'hB1, 8'hAC},
{8'h83, 8'h88, 8'h7D},
{8'h74, 8'h7C, 8'h64},
{8'hD7, 8'hDB, 8'hCA},
{8'hF3, 8'hF3, 8'hED},
{8'hF5, 8'hF1, 8'hF0},
{8'hF7, 8'hF5, 8'hF1},
{8'h91, 8'h92, 8'h83},
{8'h8A, 8'h90, 8'h72},
{8'hC4, 8'hCF, 8'hA6},
{8'hEC, 8'hF4, 8'hC3},
{8'hE1, 8'hE9, 8'hBC},
{8'hE3, 8'hEC, 8'hC4},
{8'hDA, 8'hE4, 8'hC0},
{8'hD0, 8'hDE, 8'hB6},
{8'hE1, 8'hF2, 8'hC1},
{8'hE3, 8'hF6, 8'hBD},
{8'hDC, 8'hF1, 8'hB1},
{8'hDE, 8'hF2, 8'hB6},
{8'hE0, 8'hF2, 8'hB6},
{8'hE1, 8'hF3, 8'hB6},
{8'hE5, 8'hF3, 8'hBC},
{8'hC6, 8'hD2, 8'hA8},
{8'h91, 8'h99, 8'h83},
{8'h7A, 8'h7D, 8'h79},
{8'h7D, 8'h7E, 8'h85},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'h7F, 8'h7D, 8'h81},
{8'h80, 8'h7E, 8'h82},
{8'h7A, 8'h78, 8'h7C},
{8'h96, 8'h94, 8'h97},
{8'hB0, 8'hAF, 8'hAE},
{8'h79, 8'h79, 8'h75},
{8'h9D, 8'h9C, 8'h98},
{8'hE8, 8'hE7, 8'hDF},
{8'hEA, 8'hE9, 8'hC7},
{8'hE8, 8'hE8, 8'hBB},
{8'hF1, 8'hF1, 8'hBB},
{8'hC2, 8'hC0, 8'h91},
{8'h52, 8'h4C, 8'h40},
{8'h1E, 8'h14, 8'h24},
{8'h05, 8'h00, 8'h18},
{8'h1F, 8'h18, 8'h30},
{8'hB9, 8'hB5, 8'hB9},
{8'hFF, 8'hFE, 8'hEA},
{8'hF9, 8'hFC, 8'hE6},
{8'hC8, 8'hCB, 8'hC8},
{8'h8A, 8'h8E, 8'h97},
{8'hAE, 8'hB5, 8'hBD},
{8'hA0, 8'hA4, 8'hC2},
{8'h62, 8'h60, 8'hAC},
{8'h3A, 8'h4F, 8'h98},
{8'h44, 8'h75, 8'h6D},
{8'hDF, 8'hD6, 8'h7C},
{8'hBB, 8'h9F, 8'h7F},
{8'h4F, 8'h47, 8'h5D},
{8'h66, 8'h53, 8'h41},
{8'hC6, 8'hB4, 8'h87},
{8'hDE, 8'hB8, 8'h7F},
{8'hC8, 8'h71, 8'h43},
{8'hC2, 8'h6B, 8'h47},
{8'hD0, 8'h8A, 8'h6D},
{8'hF2, 8'hDA, 8'hB8},
{8'hEB, 8'hF4, 8'hCE},
{8'hF7, 8'hFF, 8'hDE},
{8'hFA, 8'hEC, 8'hCD},
{8'hF9, 8'hC7, 8'hB4},
{8'hF7, 8'hC8, 8'hAA},
{8'hFA, 8'hCD, 8'hAA},
{8'hFB, 8'hDE, 8'hBF},
{8'hFE, 8'hF9, 8'hDA},
{8'hF7, 8'hFF, 8'hDE},
{8'hF7, 8'hFD, 8'hDA},
{8'hE0, 8'hD1, 8'hB1},
{8'hA4, 8'h7A, 8'h6A},
{8'h87, 8'h71, 8'h6F},
{8'h7D, 8'h67, 8'h58},
{8'h6A, 8'h38, 8'h1A},
{8'h97, 8'h43, 8'h1B},
{8'hCD, 8'h85, 8'h51},
{8'hF5, 8'hE3, 8'hA7},
{8'hF6, 8'hF6, 8'hC7},
{8'h93, 8'h77, 8'h5B},
{8'h8C, 8'h5B, 8'h3E},
{8'hE2, 8'hC7, 8'hA2},
{8'hD6, 8'hCA, 8'hAD},
{8'hFB, 8'hF9, 8'hEE},
{8'hF7, 8'hF3, 8'hEF},
{8'hFC, 8'hF7, 8'hF7},
{8'hFD, 8'hF9, 8'hFE},
{8'hE6, 8'hE4, 8'hE7},
{8'hA7, 8'hAE, 8'h91},
{8'hCF, 8'hD3, 8'hBE},
{8'hF2, 8'hF2, 8'hEB},
{8'hF4, 8'hF0, 8'hF0},
{8'hFF, 8'hFC, 8'hF4},
{8'hBC, 8'hBF, 8'hA7},
{8'hB5, 8'hBE, 8'h93},
{8'hE3, 8'hF0, 8'hBB},
{8'hE5, 8'hEC, 8'hC2},
{8'hE4, 8'hEA, 8'hC7},
{8'hE3, 8'hE8, 8'hCC},
{8'hF2, 8'hF8, 8'hDF},
{8'hD5, 8'hDF, 8'hC0},
{8'hD9, 8'hE8, 8'hBF},
{8'hE1, 8'hF3, 8'hBD},
{8'hDF, 8'hF5, 8'hB7},
{8'hDE, 8'hF2, 8'hB7},
{8'hE0, 8'hF3, 8'hB5},
{8'hE1, 8'hF4, 8'hB4},
{8'hE3, 8'hF3, 8'hBB},
{8'hE7, 8'hF4, 8'hC5},
{8'hE5, 8'hEF, 8'hCD},
{8'hA1, 8'hA7, 8'h98},
{8'h76, 8'h78, 8'h7A},
{8'hFF, 8'hD7, 8'h00},
{8'h7F, 8'h7D, 8'h7F},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'h7F, 8'h7D, 8'h7F},
{8'h7F, 8'h7D, 8'h7F},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'h7F, 8'h7D, 8'h81},
{8'h7E, 8'h7C, 8'h81},
{8'h85, 8'h83, 8'h87},
{8'hDA, 8'hD8, 8'hD8},
{8'hE5, 8'hE5, 8'hDF},
{8'hF2, 8'hF2, 8'hE5},
{8'hF2, 8'hF3, 8'hDF},
{8'hF3, 8'hF1, 8'hC0},
{8'hFB, 8'hF3, 8'hC0},
{8'hF3, 8'hE8, 8'h9E},
{8'hDE, 8'hD2, 8'h77},
{8'h97, 8'h89, 8'h5B},
{8'h36, 8'h28, 8'h3A},
{8'h0C, 8'h07, 8'h2C},
{8'h00, 8'h03, 8'h12},
{8'h22, 8'h1F, 8'h30},
{8'h95, 8'h97, 8'h93},
{8'hC8, 8'hD5, 8'hBF},
{8'hA0, 8'hB4, 8'hA9},
{8'h70, 8'h88, 8'hA3},
{8'h38, 8'h54, 8'h96},
{8'h22, 8'h42, 8'h97},
{8'h16, 8'h3B, 8'h92},
{8'h31, 8'h55, 8'h88},
{8'hD2, 8'hB8, 8'h77},
{8'hE4, 8'hBE, 8'h76},
{8'h39, 8'h5E, 8'h7D},
{8'h03, 8'h60, 8'hBD},
{8'h17, 8'h4B, 8'hAC},
{8'h64, 8'h4D, 8'h7B},
{8'hE7, 8'hBC, 8'h97},
{8'hBD, 8'h78, 8'h43},
{8'hC4, 8'h6A, 8'h49},
{8'hB5, 8'h53, 8'h41},
{8'hC8, 8'h87, 8'h6D},
{8'hEC, 8'hE2, 8'hB5},
{8'hF6, 8'hFF, 8'hD6},
{8'hFA, 8'hFE, 8'hDC},
{8'hFC, 8'hF4, 8'hE5},
{8'hF6, 8'hEC, 8'hEB},
{8'hF9, 8'hF6, 8'hD3},
{8'hFF, 8'hFF, 8'hD6},
{8'hFF, 8'hFF, 8'hEE},
{8'hF2, 8'hEE, 8'hDA},
{8'hD2, 8'hCA, 8'h9B},
{8'hD5, 8'hC8, 8'hA0},
{8'h96, 8'h81, 8'h7D},
{8'h83, 8'h7A, 8'h7C},
{8'h8C, 8'h75, 8'h6C},
{8'h74, 8'h30, 8'h1C},
{8'h9E, 8'h51, 8'h20},
{8'hE3, 8'hC3, 8'h76},
{8'hFF, 8'hFE, 8'hBD},
{8'hD0, 8'hB5, 8'h98},
{8'hB1, 8'h91, 8'h90},
{8'h9D, 8'h74, 8'h72},
{8'hE2, 8'hCE, 8'h98},
{8'hC7, 8'hB7, 8'h95},
{8'hFF, 8'hF8, 8'hFF},
{8'hF9, 8'hF6, 8'hEF},
{8'hF9, 8'hF8, 8'hE6},
{8'hFD, 8'hF2, 8'hF8},
{8'hFF, 8'hF6, 8'hFF},
{8'hF9, 8'hFB, 8'hDB},
{8'hE6, 8'hE8, 8'hD2},
{8'hF9, 8'hF5, 8'hF3},
{8'hFA, 8'hF4, 8'hF4},
{8'hF9, 8'hF8, 8'hE8},
{8'hD5, 8'hD9, 8'hB6},
{8'hDD, 8'hE9, 8'hB8},
{8'hE2, 8'hF2, 8'hBF},
{8'hE5, 8'hEB, 8'hD2},
{8'hEA, 8'hEC, 8'hDD},
{8'hF1, 8'hF0, 8'hE7},
{8'hF4, 8'hF1, 8'hEA},
{8'hF2, 8'hF1, 8'hE1},
{8'hE4, 8'hEC, 8'hC6},
{8'hE7, 8'hF5, 8'hB9},
{8'hDF, 8'hF4, 8'hAB},
{8'hE0, 8'hF4, 8'hC0},
{8'hE0, 8'hF6, 8'hB3},
{8'hE1, 8'hF6, 8'hB5},
{8'hE0, 8'hF1, 8'hC2},
{8'hDE, 8'hEE, 8'hBB},
{8'hE6, 8'hF7, 8'hB4},
{8'hCB, 8'hD8, 8'hAB},
{8'h7B, 8'h7F, 8'h7C},
{8'h7E, 8'h7D, 8'h7B},
{8'h7F, 8'h7E, 8'h7C},
{8'h7F, 8'h7D, 8'h7E},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'h7F, 8'h7D, 8'h7E},
{8'h7F, 8'h7E, 8'h7C},
{8'h7F, 8'h7E, 8'h7B},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'h7F, 8'h7D, 8'h7F},
{8'hFF, 8'hD7, 8'h00},
{8'h7F, 8'h7D, 8'h82},
{8'h7C, 8'h7A, 8'h7E},
{8'h98, 8'h97, 8'h97},
{8'hED, 8'hED, 8'hE7},
{8'hFA, 8'hFB, 8'hEE},
{8'hFA, 8'hFB, 8'hEB},
{8'hF8, 8'hF4, 8'hE0},
{8'hF8, 8'hF1, 8'hD3},
{8'hF9, 8'hEE, 8'hC0},
{8'hF9, 8'hEE, 8'hB4},
{8'hFD, 8'hF5, 8'hC8},
{8'hE8, 8'hE2, 8'hD5},
{8'hB8, 8'hBA, 8'hC0},
{8'hB7, 8'hBE, 8'hC0},
{8'hC1, 8'hCA, 8'hB0},
{8'hA1, 8'hAF, 8'hA0},
{8'h61, 8'h6E, 8'h83},
{8'h25, 8'h31, 8'h75},
{8'h09, 8'h17, 8'h7A},
{8'h06, 8'h12, 8'h6C},
{8'h00, 8'h19, 8'h46},
{8'h00, 8'h18, 8'h24},
{8'h06, 8'h0D, 8'h2C},
{8'h28, 8'h21, 8'h17},
{8'h2F, 8'h1F, 8'h19},
{8'h24, 8'h2B, 8'h5C},
{8'h1F, 8'h55, 8'hAE},
{8'h18, 8'h59, 8'hC5},
{8'h29, 8'h42, 8'h76},
{8'h87, 8'h75, 8'h43},
{8'hC7, 8'h93, 8'h58},
{8'hA9, 8'h61, 8'h38},
{8'hAC, 8'h4B, 8'h34},
{8'hB6, 8'h48, 8'h39},
{8'hE4, 8'h8B, 8'h78},
{8'hFF, 8'hE4, 8'hC7},
{8'hFF, 8'hFF, 8'hDE},
{8'hF1, 8'hFD, 8'hDF},
{8'hFB, 8'hFE, 8'hE0},
{8'hFF, 8'hFF, 8'hDA},
{8'hFA, 8'hED, 8'hD4},
{8'hB9, 8'h98, 8'hA3},
{8'h68, 8'h47, 8'h4E},
{8'hC9, 8'hB8, 8'h99},
{8'hFE, 8'hFF, 8'hCD},
{8'hB4, 8'hC1, 8'h9B},
{8'h69, 8'h7B, 8'h8E},
{8'h74, 8'h86, 8'h8B},
{8'h76, 8'h34, 8'h34},
{8'hCB, 8'h7B, 8'h5F},
{8'hFC, 8'hFC, 8'hB8},
{8'hF4, 8'hF7, 8'hB4},
{8'hAA, 8'h78, 8'h56},
{8'hEB, 8'hD2, 8'hBD},
{8'hBF, 8'hAA, 8'h8A},
{8'hE3, 8'hDB, 8'h9A},
{8'hAC, 8'h9F, 8'h85},
{8'hDE, 8'hD0, 8'hE6},
{8'hFA, 8'hF6, 8'hFA},
{8'hF5, 8'hF5, 8'hE7},
{8'hFB, 8'hF9, 8'hF1},
{8'hF9, 8'hF8, 8'hEB},
{8'hFE, 8'hFB, 8'hFF},
{8'hFA, 8'hF3, 8'hFF},
{8'hF9, 8'hF1, 8'hFD},
{8'hFD, 8'hF6, 8'hF5},
{8'hF8, 8'hF4, 8'hE9},
{8'hEF, 8'hEE, 8'hE5},
{8'hE8, 8'hEB, 8'hEC},
{8'hEA, 8'hEF, 8'hF6},
{8'hF3, 8'hF7, 8'hEC},
{8'hF2, 8'hF2, 8'hEC},
{8'hEF, 8'hEC, 8'hEE},
{8'hEE, 8'hE9, 8'hEB},
{8'hF2, 8'hF0, 8'hE8},
{8'hE4, 8'hE9, 8'hCE},
{8'hDF, 8'hEC, 8'hBC},
{8'hDD, 8'hEF, 8'hB3},
{8'hE1, 8'hF5, 8'hBF},
{8'hE1, 8'hF7, 8'hB2},
{8'hE1, 8'hF6, 8'hB4},
{8'hE1, 8'hF1, 8'hC3},
{8'hE1, 8'hF0, 8'hBE},
{8'hE7, 8'hF9, 8'hB5},
{8'hE9, 8'hF6, 8'hC8},
{8'h9B, 8'h9F, 8'h9B},
{8'h7C, 8'h7A, 8'h7D},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'h7F, 8'h7D, 8'h7E},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'h7F, 8'h7D, 8'h7E},
{8'hFF, 8'hD7, 8'h00},
{8'h7F, 8'h7D, 8'h82},
{8'h7F, 8'h7D, 8'h82},
{8'h7A, 8'h78, 8'h7B},
{8'h8C, 8'h8B, 8'h88},
{8'hC4, 8'hC4, 8'hBB},
{8'hD8, 8'hD8, 8'hCD},
{8'hF6, 8'hF3, 8'hF4},
{8'hFA, 8'hF5, 8'hE9},
{8'hFE, 8'hF5, 8'hE3},
{8'hFE, 8'hF5, 8'hE3},
{8'hF6, 8'hF0, 8'hD1},
{8'hF8, 8'hFA, 8'hD1},
{8'hF8, 8'hFD, 8'hEC},
{8'h99, 8'hA2, 8'hB4},
{8'h45, 8'h5D, 8'h92},
{8'h1A, 8'h36, 8'h73},
{8'h15, 8'h2E, 8'h7D},
{8'h19, 8'h31, 8'h98},
{8'h1B, 8'h36, 8'hAF},
{8'h1C, 8'h39, 8'hAE},
{8'h17, 8'h3E, 8'h9A},
{8'h19, 8'h3A, 8'h80},
{8'h1B, 8'h1E, 8'h5D},
{8'h01, 8'h15, 8'h4C},
{8'h00, 8'h02, 8'h34},
{8'h07, 8'h00, 8'h26},
{8'h16, 8'h22, 8'h59},
{8'h13, 8'h54, 8'hB5},
{8'h12, 8'h51, 8'h9A},
{8'h33, 8'h41, 8'h33},
{8'hAE, 8'h76, 8'h47},
{8'h9D, 8'h5C, 8'h32},
{8'h8A, 8'h38, 8'h18},
{8'h95, 8'h29, 8'h17},
{8'hAA, 8'h30, 8'h27},
{8'hC8, 8'h70, 8'h64},
{8'hF2, 8'hD5, 8'hBB},
{8'hFF, 8'hFF, 8'hE1},
{8'hFC, 8'hF7, 8'hCF},
{8'hC3, 8'hAA, 8'h86},
{8'h5A, 8'h3B, 8'h31},
{8'h20, 8'h00, 8'h12},
{8'h18, 8'h04, 8'h0F},
{8'hA0, 8'h98, 8'h81},
{8'hF5, 8'hFD, 8'hC5},
{8'hEA, 8'hF5, 8'hBE},
{8'h9B, 8'h8F, 8'h89},
{8'h72, 8'h5F, 8'h50},
{8'h9E, 8'h78, 8'h5B},
{8'hFF, 8'hE9, 8'hBF},
{8'hFF, 8'hF9, 8'hC9},
{8'hB1, 8'hA7, 8'h7F},
{8'hA5, 8'h9E, 8'h87},
{8'hFF, 8'hFF, 8'hF6},
{8'hE7, 8'hDE, 8'hBC},
{8'hE1, 8'hDA, 8'h99},
{8'hA0, 8'h95, 8'h73},
{8'h93, 8'h85, 8'h88},
{8'hE6, 8'hE0, 8'hCE},
{8'hFA, 8'hF9, 8'hE1},
{8'hFA, 8'hFB, 8'hF2},
{8'hF4, 8'hF7, 8'hE7},
{8'hF9, 8'hF6, 8'hF3},
{8'hFB, 8'hF6, 8'hF2},
{8'hF9, 8'hF2, 8'hE7},
{8'hFC, 8'hF5, 8'hE2},
{8'hF9, 8'hF4, 8'hE1},
{8'hF6, 8'hF5, 8'hE6},
{8'hF5, 8'hF6, 8'hEF},
{8'hF1, 8'hF5, 8'hEF},
{8'hF3, 8'hF5, 8'hEF},
{8'hF5, 8'hF3, 8'hF2},
{8'hF7, 8'hF1, 8'hF7},
{8'hF8, 8'hF1, 8'hF6},
{8'hF1, 8'hED, 8'hEA},
{8'hD8, 8'hDB, 8'hC7},
{8'hE2, 8'hED, 8'hC6},
{8'hE2, 8'hF2, 8'hBF},
{8'hE2, 8'hF4, 8'hBE},
{8'hE1, 8'hF7, 8'hB0},
{8'hE2, 8'hF5, 8'hB4},
{8'hE3, 8'hF2, 8'hC5},
{8'hE1, 8'hEF, 8'hBE},
{8'hE8, 8'hF7, 8'hB6},
{8'hD6, 8'hE2, 8'hB3},
{8'hA8, 8'hAC, 8'hA6},
{8'h7C, 8'h79, 8'h81},
{8'h7F, 8'h7C, 8'h82},
{8'h7F, 8'h7D, 8'h82},
{8'h7F, 8'h7D, 8'h82},
{8'h7F, 8'h7D, 8'h81},
{8'h7F, 8'h7D, 8'h82},
{8'h7F, 8'h7C, 8'h83},
{8'h7F, 8'h7C, 8'h83},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'h7F, 8'h7D, 8'h7D},
{8'h7F, 8'h7D, 8'h7F},
{8'h7F, 8'h7D, 8'h82},
{8'h7F, 8'h7D, 8'h83},
{8'h84, 8'h82, 8'h86},
{8'h7C, 8'h7A, 8'h7A},
{8'h76, 8'h76, 8'h71},
{8'h89, 8'h89, 8'h81},
{8'hF1, 8'hF1, 8'hF0},
{8'hFC, 8'hFC, 8'hED},
{8'hFB, 8'hF8, 8'hEF},
{8'hF7, 8'hF0, 8'hF6},
{8'hF4, 8'hF1, 8'hE2},
{8'hFE, 8'hFF, 8'hD6},
{8'hE3, 8'hEA, 8'hD8},
{8'h34, 8'h39, 8'h6B},
{8'h14, 8'h43, 8'hBA},
{8'h1A, 8'h4F, 8'hBE},
{8'h1F, 8'h55, 8'hB5},
{8'h1A, 8'h52, 8'hAB},
{8'h1E, 8'h55, 8'hB1},
{8'h1E, 8'h54, 8'hBA},
{8'h1B, 8'h50, 8'hC2},
{8'h1F, 8'h50, 8'hC8},
{8'h31, 8'h4C, 8'hBA},
{8'h18, 8'h53, 8'hBD},
{8'h08, 8'h38, 8'h83},
{8'h08, 8'h0B, 8'h26},
{8'h02, 8'h00, 8'h15},
{8'h03, 8'h20, 8'h65},
{8'h1E, 8'h55, 8'hAB},
{8'h18, 8'h2B, 8'h63},
{8'h82, 8'h41, 8'h2E},
{8'hA1, 8'h5F, 8'h3E},
{8'h6D, 8'h2E, 8'h0C},
{8'h5B, 8'h1E, 8'h04},
{8'h62, 8'h25, 8'h11},
{8'h67, 8'h27, 8'h1A},
{8'h7A, 8'h39, 8'h29},
{8'hBF, 8'h85, 8'h71},
{8'h99, 8'h5B, 8'h48},
{8'h51, 8'h1D, 8'h0E},
{8'h16, 8'h00, 8'h00},
{8'h1B, 8'h19, 8'h17},
{8'h97, 8'hA2, 8'h98},
{8'hF1, 8'hFA, 8'hE1},
{8'hF2, 8'hF3, 8'hCA},
{8'hFB, 8'hF3, 8'hC8},
{8'hCA, 8'hA3, 8'h8C},
{8'hAF, 8'hA1, 8'h74},
{8'hF2, 8'hF2, 8'hB7},
{8'hEE, 8'hDE, 8'hA4},
{8'hE3, 8'hB1, 8'h8B},
{8'h9F, 8'h57, 8'h43},
{8'hCD, 8'hA1, 8'h8C},
{8'hDF, 8'hDD, 8'hC2},
{8'hF3, 8'hE9, 8'hD1},
{8'hF1, 8'hE7, 8'hB1},
{8'hB1, 8'hA5, 8'h78},
{8'hDA, 8'hD0, 8'hAE},
{8'hDC, 8'hD9, 8'hA4},
{8'hDE, 8'hDE, 8'hBD},
{8'hFE, 8'hFD, 8'hFF},
{8'hF8, 8'hF9, 8'hF4},
{8'hF8, 8'hF6, 8'hE0},
{8'hF8, 8'hF4, 8'hDB},
{8'hFE, 8'hFA, 8'hE2},
{8'hFF, 8'hF7, 8'hE9},
{8'hFA, 8'hF0, 8'hEB},
{8'hF4, 8'hEF, 8'hEA},
{8'hFD, 8'hFD, 8'hEE},
{8'hF4, 8'hF9, 8'hE0},
{8'hF9, 8'hFA, 8'hED},
{8'hF8, 8'hF6, 8'hEF},
{8'hF5, 8'hF0, 8'hED},
{8'hF5, 8'hEF, 8'hEB},
{8'hE2, 8'hDE, 8'hD2},
{8'hE4, 8'hE6, 8'hCC},
{8'hE9, 8'hF2, 8'hC8},
{8'hE3, 8'hF1, 8'hBE},
{8'hE1, 8'hF3, 8'hBC},
{8'hE2, 8'hF7, 8'hB1},
{8'hE2, 8'hF4, 8'hB6},
{8'hE3, 8'hF0, 8'hC9},
{8'hE4, 8'hEF, 8'hC4},
{8'hEC, 8'hF9, 8'hBB},
{8'hBD, 8'hC6, 8'h98},
{8'h7A, 8'h7D, 8'h77},
{8'h7E, 8'h7B, 8'h86},
{8'h7D, 8'h7A, 8'h82},
{8'h7F, 8'h7D, 8'h82},
{8'h7F, 8'h7D, 8'h7F},
{8'h82, 8'h80, 8'h82},
{8'h7F, 8'h7D, 8'h82},
{8'h80, 8'h7D, 8'h85},
{8'h7F, 8'h7C, 8'h85},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'h7F, 8'h7E, 8'h7C},
{8'h7F, 8'h7D, 8'h7F},
{8'h7F, 8'h7D, 8'h82},
{8'h7E, 8'h7B, 8'h82},
{8'h7B, 8'h79, 8'h7F},
{8'h81, 8'h7F, 8'h82},
{8'h7F, 8'h7E, 8'h7B},
{8'hA3, 8'hA3, 8'h9D},
{8'hF1, 8'hF3, 8'hE3},
{8'hFD, 8'hFE, 8'hE5},
{8'hF0, 8'hF0, 8'hE3},
{8'hF5, 8'hF2, 8'hF8},
{8'hF9, 8'hF8, 8'hF2},
{8'hFA, 8'hFD, 8'hE2},
{8'hDE, 8'hE0, 8'hDE},
{8'h24, 8'h26, 8'h5D},
{8'h0F, 8'h57, 8'hAD},
{8'h0A, 8'h57, 8'hB1},
{8'h0C, 8'h57, 8'hB3},
{8'h0F, 8'h59, 8'hB0},
{8'h0F, 8'h5A, 8'hA8},
{8'h0F, 8'h58, 8'hA3},
{8'h10, 8'h58, 8'hA7},
{8'h13, 8'h59, 8'hAE},
{8'h16, 8'h58, 8'hC1},
{8'h08, 8'h52, 8'hC1},
{8'h16, 8'h5C, 8'hB4},
{8'h16, 8'h3D, 8'h75},
{8'h03, 8'h08, 8'h36},
{8'h01, 8'h00, 8'h2F},
{8'h10, 8'h22, 8'h64},
{8'h16, 8'h32, 8'h85},
{8'h3B, 8'h1D, 8'h1D},
{8'h92, 8'h5E, 8'h4A},
{8'h67, 8'h31, 8'h15},
{8'h36, 8'h17, 8'h02},
{8'h1F, 8'h1A, 8'h09},
{8'h26, 8'h1C, 8'h11},
{8'h4B, 8'h16, 8'h0F},
{8'h6C, 8'h0D, 8'h07},
{8'h5E, 8'h16, 8'h17},
{8'h49, 8'h15, 8'h1A},
{8'h78, 8'h61, 8'h5C},
{8'hD4, 8'hD7, 8'hC1},
{8'hEF, 8'hFA, 8'hE0},
{8'hF4, 8'hFC, 8'hE9},
{8'hF7, 8'hF8, 8'hE5},
{8'hF2, 8'hEB, 8'hD2},
{8'hEC, 8'hD3, 8'hB7},
{8'hE0, 8'hF2, 8'hB9},
{8'hC0, 8'hB5, 8'h73},
{8'hDD, 8'hAA, 8'h79},
{8'h98, 8'h68, 8'h40},
{8'hA7, 8'h4A, 8'h34},
{8'hBE, 8'h46, 8'h2C},
{8'h85, 8'h50, 8'h1F},
{8'h8D, 8'h75, 8'h51},
{8'hD1, 8'hC2, 8'h91},
{8'hB4, 8'hA6, 8'h90},
{8'hBB, 8'hB8, 8'hAA},
{8'hB6, 8'hBA, 8'h9A},
{8'hAB, 8'hAD, 8'hA5},
{8'hBC, 8'hBD, 8'hCB},
{8'hF4, 8'hF6, 8'hEC},
{8'hFA, 8'hF3, 8'hF1},
{8'hF9, 8'hF2, 8'hDF},
{8'hF9, 8'hF2, 8'hCE},
{8'hF7, 8'hEE, 8'hCF},
{8'hF9, 8'hEE, 8'hE4},
{8'hF1, 8'hE7, 8'hED},
{8'hF0, 8'hEB, 8'hF1},
{8'hF9, 8'hF7, 8'hF5},
{8'hF6, 8'hF8, 8'hE3},
{8'hE3, 8'hE1, 8'hCF},
{8'hEA, 8'hE5, 8'hD5},
{8'hE3, 8'hDD, 8'hCD},
{8'hF3, 8'hF1, 8'hD9},
{8'hF0, 8'hF2, 8'hCE},
{8'hE4, 8'hED, 8'hBC},
{8'hDF, 8'hED, 8'hB5},
{8'hE6, 8'hF6, 8'hC1},
{8'hE4, 8'hF6, 8'hB5},
{8'hDC, 8'hEB, 8'hB4},
{8'hE2, 8'hEC, 8'hCC},
{8'hE3, 8'hEC, 8'hC9},
{8'hE6, 8'hF1, 8'hB9},
{8'hE7, 8'hEE, 8'hC5},
{8'h97, 8'h99, 8'h95},
{8'h7F, 8'h7C, 8'h87},
{8'h81, 8'h7E, 8'h85},
{8'h7E, 8'h7C, 8'h7E},
{8'h7C, 8'h7B, 8'h78},
{8'h81, 8'h80, 8'h7D},
{8'h80, 8'h7E, 8'h80},
{8'h7E, 8'h7B, 8'h83},
{8'h7E, 8'h7B, 8'h86},
{8'h7F, 8'h7D, 8'h81},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'h7F, 8'h7E, 8'h7B},
{8'h7F, 8'h7E, 8'h7E},
{8'h7F, 8'h7D, 8'h81},
{8'h7F, 8'h7C, 8'h84},
{8'h81, 8'h7E, 8'h86},
{8'h7D, 8'h7A, 8'h80},
{8'h7D, 8'h7C, 8'h7D},
{8'h7A, 8'h78, 8'h75},
{8'hAF, 8'hB2, 8'h99},
{8'hD9, 8'hDC, 8'hC0},
{8'hDD, 8'hDF, 8'hCB},
{8'hF3, 8'hF3, 8'hEA},
{8'hFB, 8'hFA, 8'hF5},
{8'hFE, 8'hFD, 8'hFB},
{8'hEC, 8'hE8, 8'hEE},
{8'h1D, 8'h1C, 8'h3D},
{8'h0C, 8'h50, 8'hA9},
{8'h0F, 8'h58, 8'hBF},
{8'h0D, 8'h52, 8'hC0},
{8'h10, 8'h56, 8'hBD},
{8'h0F, 8'h56, 8'hAD},
{8'h13, 8'h5A, 8'hAB},
{8'h14, 8'h59, 8'hB3},
{8'h12, 8'h55, 8'hB8},
{8'h08, 8'h57, 8'hA2},
{8'h13, 8'h58, 8'hB7},
{8'h16, 8'h5A, 8'hBB},
{8'h19, 8'h57, 8'hB6},
{8'h12, 8'h2A, 8'h83},
{8'h07, 8'h00, 8'h2B},
{8'h04, 8'h02, 8'h1C},
{8'h1C, 8'h2F, 8'h6E},
{8'h07, 8'h0A, 8'h16},
{8'h5D, 8'h45, 8'h3F},
{8'h57, 8'h2B, 8'h21},
{8'h34, 8'h18, 8'h10},
{8'h00, 8'h01, 8'h03},
{8'h00, 8'h02, 8'h0A},
{8'h18, 8'h02, 8'h04},
{8'h49, 8'h11, 8'h09},
{8'h3B, 8'h14, 8'h0F},
{8'h29, 8'h08, 8'h12},
{8'hCD, 8'hB5, 8'hBE},
{8'hFF, 8'hFF, 8'hF3},
{8'hFF, 8'hFD, 8'hE8},
{8'hFE, 8'hFD, 8'hF9},
{8'hCC, 8'hD0, 8'hCB},
{8'hC3, 8'hCA, 8'hAE},
{8'hF2, 8'hE1, 8'hA6},
{8'hB1, 8'h90, 8'h4A},
{8'hC4, 8'h83, 8'h48},
{8'hAF, 8'h6C, 8'h4B},
{8'h4F, 8'h32, 8'h26},
{8'h2B, 8'h0E, 8'h10},
{8'h76, 8'h3C, 8'h38},
{8'hDD, 8'hA7, 8'h8D},
{8'hC4, 8'hA8, 8'h6F},
{8'h85, 8'h78, 8'h56},
{8'h31, 8'h2C, 8'h45},
{8'h01, 8'h09, 8'h39},
{8'h04, 8'h18, 8'h3A},
{8'h13, 8'h27, 8'h57},
{8'h2F, 8'h3E, 8'h66},
{8'hBC, 8'hCB, 8'hBC},
{8'hF9, 8'hF1, 8'hEC},
{8'hF5, 8'hEF, 8'hC2},
{8'hE9, 8'hE9, 8'h8A},
{8'hE5, 8'hE4, 8'h7C},
{8'hF0, 8'hEC, 8'hA3},
{8'hF2, 8'hEA, 8'hCC},
{8'hF3, 8'hEC, 8'hE8},
{8'hF4, 8'hF0, 8'hF0},
{8'hED, 8'hEC, 8'hD8},
{8'hD8, 8'hD6, 8'hC1},
{8'hE9, 8'hE3, 8'hD0},
{8'hE7, 8'hE1, 8'hCC},
{8'hFD, 8'hFA, 8'hDF},
{8'hF2, 8'hF4, 8'hCE},
{8'hE6, 8'hED, 8'hBE},
{8'hE1, 8'hED, 8'hB9},
{8'hE2, 8'hF0, 8'hC0},
{8'hE6, 8'hF5, 8'hBA},
{8'hCE, 8'hDA, 8'hAC},
{8'h89, 8'h91, 8'h7D},
{8'hB5, 8'hBA, 8'hA1},
{8'hE9, 8'hF2, 8'hC3},
{8'hEA, 8'hF0, 8'hCC},
{8'h9C, 8'h9B, 8'h9C},
{8'h78, 8'h75, 8'h7F},
{8'hFF, 8'hD7, 8'h00},
{8'h79, 8'h78, 8'h74},
{8'h85, 8'h84, 8'h7A},
{8'h82, 8'h82, 8'h77},
{8'h7D, 8'h7C, 8'h77},
{8'h79, 8'h77, 8'h7B},
{8'h82, 8'h7F, 8'h88},
{8'h80, 8'h7E, 8'h81},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'h7F, 8'h7E, 8'h7A},
{8'h7F, 8'h7E, 8'h7D},
{8'h7F, 8'h7D, 8'h81},
{8'h7F, 8'h7B, 8'h84},
{8'h7E, 8'h7A, 8'h84},
{8'h81, 8'h7E, 8'h85},
{8'h7D, 8'h7B, 8'h80},
{8'h79, 8'h77, 8'h78},
{8'h84, 8'h83, 8'h74},
{8'h75, 8'h73, 8'h68},
{8'hA9, 8'hAA, 8'h97},
{8'hD5, 8'hD8, 8'hBB},
{8'hE8, 8'hE8, 8'hDC},
{8'hFF, 8'hFC, 8'hFF},
{8'hF8, 8'hF1, 8'hF5},
{8'h37, 8'h34, 8'h34},
{8'h01, 8'h30, 8'h81},
{8'h1E, 8'h54, 8'hBA},
{8'h1B, 8'h4F, 8'hC1},
{8'h1B, 8'h4F, 8'hBA},
{8'h1D, 8'h54, 8'hAC},
{8'h18, 8'h50, 8'h9F},
{8'h18, 8'h4D, 8'hAA},
{8'h1C, 8'h4E, 8'hB9},
{8'h1D, 8'h51, 8'h94},
{8'h20, 8'h50, 8'hB3},
{8'h16, 8'h56, 8'hB5},
{8'h11, 8'h5A, 8'hB0},
{8'h1C, 8'h4A, 8'h9F},
{8'h05, 8'h0C, 8'h32},
{8'h04, 8'h02, 8'h0E},
{8'h0F, 8'h12, 8'h44},
{8'h10, 8'h0B, 8'h33},
{8'h26, 8'h1D, 8'h27},
{8'h3B, 8'h2B, 8'h26},
{8'h29, 8'h1C, 8'h1A},
{8'h06, 8'h00, 8'h15},
{8'h06, 8'h00, 8'h22},
{8'h07, 8'h00, 8'h0E},
{8'h26, 8'h19, 8'h0D},
{8'h3C, 8'h1E, 8'h05},
{8'h16, 8'h02, 8'h07},
{8'h53, 8'h47, 8'h5D},
{8'h94, 8'h96, 8'h97},
{8'hB4, 8'hB8, 8'hB5},
{8'h95, 8'h93, 8'h9F},
{8'h49, 8'h45, 8'h44},
{8'hE0, 8'hDC, 8'hB4},
{8'hC4, 8'h97, 8'h68},
{8'h94, 8'h51, 8'h24},
{8'hAD, 8'h5F, 8'h3D},
{8'h56, 8'h26, 8'h20},
{8'h24, 8'h22, 8'h40},
{8'h08, 8'h1E, 8'h4A},
{8'h10, 8'h1D, 8'h39},
{8'h2B, 8'h1F, 8'h23},
{8'h5E, 8'h41, 8'h27},
{8'h33, 8'h28, 8'h28},
{8'h14, 8'h23, 8'h64},
{8'h15, 8'h46, 8'h9B},
{8'h1A, 8'h5C, 8'hA5},
{8'h1C, 8'h54, 8'hB5},
{8'h22, 8'h48, 8'hA1},
{8'h5A, 8'h78, 8'h8B},
{8'hFD, 8'hF7, 8'hE6},
{8'hEF, 8'hEA, 8'hA9},
{8'hD4, 8'hD6, 8'h62},
{8'hDC, 8'hDD, 8'h66},
{8'hE6, 8'hE1, 8'h92},
{8'hF4, 8'hEC, 8'hCA},
{8'hF9, 8'hF3, 8'hE5},
{8'hF2, 8'hEE, 8'hE1},
{8'hF5, 8'hF3, 8'hE6},
{8'hF3, 8'hEE, 8'hE2},
{8'hD8, 8'hD0, 8'hC4},
{8'hF4, 8'hED, 8'hDF},
{8'hFD, 8'hFB, 8'hE8},
{8'hEB, 8'hEA, 8'hCE},
{8'hDE, 8'hE3, 8'hBF},
{8'hE2, 8'hEB, 8'hC3},
{8'hE4, 8'hF1, 8'hC6},
{8'hE4, 8'hF1, 8'hBC},
{8'hD9, 8'hE4, 8'hBD},
{8'h80, 8'h84, 8'h79},
{8'h97, 8'h9B, 8'h8B},
{8'hEC, 8'hF2, 8'hCA},
{8'hB0, 8'hB4, 8'h96},
{8'h7D, 8'h7A, 8'h80},
{8'h7B, 8'h77, 8'h80},
{8'h76, 8'h75, 8'h75},
{8'h91, 8'h90, 8'h87},
{8'hD3, 8'hD4, 8'hC3},
{8'h96, 8'h97, 8'h85},
{8'h7A, 8'h7A, 8'h6F},
{8'h7C, 8'h7B, 8'h7B},
{8'h81, 8'h7E, 8'h85},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'h7F, 8'h7D, 8'h7F},
{8'h80, 8'h7E, 8'h80},
{8'h7F, 8'h7D, 8'h7E},
{8'h7F, 8'h7D, 8'h7E},
{8'h81, 8'h7C, 8'h7F},
{8'h81, 8'h7C, 8'h7F},
{8'h80, 8'h7D, 8'h81},
{8'h7B, 8'h7C, 8'h82},
{8'h7B, 8'h7F, 8'h85},
{8'h78, 8'h7C, 8'h80},
{8'h96, 8'h97, 8'h95},
{8'hCF, 8'hCC, 8'hC5},
{8'hED, 8'hEA, 8'hDC},
{8'hBD, 8'hBC, 8'hB3},
{8'h7E, 8'h80, 8'h6C},
{8'hD1, 8'hD3, 8'hB1},
{8'hF8, 8'hF0, 8'hE5},
{8'hED, 8'hDB, 8'hE6},
{8'hE4, 8'hD9, 8'hD7},
{8'h7C, 8'h7B, 8'h65},
{8'h12, 8'h33, 8'h41},
{8'h24, 8'h4B, 8'h80},
{8'h2E, 8'h4D, 8'hA2},
{8'h18, 8'h34, 8'h89},
{8'h0E, 8'h21, 8'h67},
{8'h0E, 8'h28, 8'h65},
{8'h08, 8'h35, 8'h77},
{8'h13, 8'h4B, 8'h8F},
{8'h24, 8'h42, 8'h93},
{8'h11, 8'h2E, 8'h96},
{8'h04, 8'h34, 8'h88},
{8'h11, 8'h58, 8'h97},
{8'h21, 8'h59, 8'h9D},
{8'h0C, 8'h23, 8'h4C},
{8'h00, 8'h01, 8'h14},
{8'h07, 8'h01, 8'h2C},
{8'h19, 8'h01, 8'h35},
{8'h09, 8'h02, 8'h1E},
{8'h15, 8'h20, 8'h2F},
{8'h17, 8'h2D, 8'h48},
{8'h05, 8'h10, 8'h38},
{8'h09, 8'h01, 8'h27},
{8'h04, 8'h00, 8'h0C},
{8'h12, 8'h17, 8'h08},
{8'h45, 8'h21, 8'h00},
{8'h22, 8'h06, 8'h0A},
{8'h00, 8'h00, 8'h19},
{8'h00, 8'h00, 8'h1B},
{8'h03, 8'h1A, 8'h34},
{8'h18, 8'h25, 8'h44},
{8'h8B, 8'h7A, 8'h7E},
{8'hE2, 8'hBE, 8'h9B},
{8'h60, 8'h2F, 8'h30},
{8'h27, 8'h15, 8'h0C},
{8'h5E, 8'h3A, 8'h34},
{8'h21, 8'h06, 8'h1E},
{8'h23, 8'h39, 8'h68},
{8'h06, 8'h1D, 8'h4D},
{8'h03, 8'h02, 8'h21},
{8'h04, 8'h16, 8'h19},
{8'h30, 8'h2A, 8'h3E},
{8'h19, 8'h20, 8'h4C},
{8'h23, 8'h4A, 8'h9C},
{8'h18, 8'h5C, 8'hB3},
{8'h0C, 8'h5D, 8'hA9},
{8'h0E, 8'h52, 8'hBD},
{8'h24, 8'h55, 8'hC5},
{8'h1F, 8'h3B, 8'h75},
{8'hDC, 8'hD1, 8'hC7},
{8'hF8, 8'hEE, 8'hC4},
{8'hE8, 8'hE0, 8'h9C},
{8'hF4, 8'hEB, 8'hAF},
{8'hFF, 8'hF6, 8'hDD},
{8'hFD, 8'hF0, 8'hF2},
{8'hFA, 8'hF0, 8'hF7},
{8'hFA, 8'hF4, 8'hF2},
{8'hF9, 8'hF6, 8'hF4},
{8'hFD, 8'hF8, 8'hF5},
{8'hF0, 8'hE9, 8'hE6},
{8'hEB, 8'hE4, 8'hDD},
{8'hF5, 8'hEE, 8'hE3},
{8'hF7, 8'hF5, 8'hE3},
{8'hF1, 8'hF3, 8'hDC},
{8'hE8, 8'hEC, 8'hD2},
{8'hE5, 8'hED, 8'hCB},
{8'hD0, 8'hD9, 8'hAF},
{8'hAF, 8'hB7, 8'h97},
{8'hC0, 8'hC3, 8'hB8},
{8'h7A, 8'h7C, 8'h6F},
{8'h95, 8'h9A, 8'h7C},
{8'h7E, 8'h81, 8'h6C},
{8'h7D, 8'h7C, 8'h83},
{8'h7C, 8'h7D, 8'h7B},
{8'h8D, 8'h90, 8'h84},
{8'hE0, 8'hE3, 8'hD1},
{8'hC2, 8'hC5, 8'hB3},
{8'h7D, 8'h7E, 8'h72},
{8'h7F, 8'h80, 8'h7A},
{8'h7E, 8'h7E, 8'h78},
{8'h85, 8'h86, 8'h7E},
{8'h7F, 8'h7E, 8'h7F},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'h7F, 8'h7D, 8'h82},
{8'h7F, 8'h7D, 8'h81},
{8'hFF, 8'hD7, 8'h00},
{8'h7F, 8'h7D, 8'h7F},
{8'h7E, 8'h7D, 8'h7C},
{8'h82, 8'h81, 8'h7F},
{8'h85, 8'h84, 8'h80},
{8'h7C, 8'h7B, 8'h78},
{8'h85, 8'h76, 8'h8A},
{8'h84, 8'h76, 8'h82},
{8'h7B, 8'h76, 8'h77},
{8'h79, 8'h83, 8'h7F},
{8'h6F, 8'h84, 8'h80},
{8'h70, 8'h82, 8'h77},
{8'hB3, 8'hB2, 8'h9B},
{8'hE7, 8'hD5, 8'hB2},
{8'hE5, 8'hDE, 8'hB7},
{8'hDB, 8'hE3, 8'hBD},
{8'hB7, 8'hC8, 8'hA7},
{8'hE4, 8'hE7, 8'hD2},
{8'hEB, 8'hD6, 8'hCC},
{8'hFA, 8'hE5, 8'hDD},
{8'hFD, 8'hF7, 8'hE6},
{8'hFC, 8'hFF, 8'hE6},
{8'hD0, 8'hDF, 8'hD2},
{8'h7D, 8'h88, 8'h9C},
{8'h1C, 8'h20, 8'h53},
{8'h0D, 8'h17, 8'h4F},
{8'h16, 8'h33, 8'h71},
{8'h14, 8'h42, 8'h8F},
{8'h08, 8'h46, 8'h99},
{8'h03, 8'h42, 8'h90},
{8'h1F, 8'h48, 8'hA2},
{8'h22, 8'h55, 8'hA4},
{8'h13, 8'h4A, 8'h92},
{8'h0E, 8'h47, 8'h9A},
{8'h22, 8'h52, 8'hAF},
{8'h14, 8'h2A, 8'h79},
{8'h00, 8'h01, 8'h2A},
{8'h06, 8'h03, 8'h0A},
{8'h09, 8'h01, 8'h12},
{8'h0A, 8'h00, 8'h1B},
{8'h02, 8'h09, 8'h46},
{8'h12, 8'h48, 8'hB0},
{8'h0F, 8'h50, 8'hB7},
{8'h18, 8'h3B, 8'h7B},
{8'h10, 8'h27, 8'h46},
{8'h08, 8'h1D, 8'h39},
{8'h19, 8'h0E, 8'h38},
{8'h31, 8'h26, 8'h09},
{8'h4B, 8'h4D, 8'h31},
{8'h25, 8'h39, 8'h87},
{8'h1E, 8'h4F, 8'hCB},
{8'h20, 8'h56, 8'h8D},
{8'h92, 8'h9E, 8'h9F},
{8'h71, 8'h51, 8'h5E},
{8'h00, 8'h00, 8'h03},
{8'h14, 8'h17, 8'h0D},
{8'h1E, 8'h1D, 8'h22},
{8'h0B, 8'h06, 8'h37},
{8'h38, 8'h34, 8'h76},
{8'h02, 8'h06, 8'h30},
{8'h03, 8'h0F, 8'h33},
{8'h25, 8'h43, 8'h7D},
{8'h10, 8'h46, 8'h9A},
{8'h15, 8'h4E, 8'hA4},
{8'h1C, 8'h59, 8'hAF},
{8'h18, 8'h56, 8'hAD},
{8'h1C, 8'h56, 8'hAD},
{8'h1A, 8'h51, 8'hA4},
{8'h1E, 8'h53, 8'hA3},
{8'h0F, 8'h3A, 8'h82},
{8'h96, 8'h91, 8'h87},
{8'hFF, 8'hFB, 8'hE3},
{8'hF2, 8'hEB, 8'hCD},
{8'hEC, 8'hE9, 8'hC8},
{8'hEE, 8'hED, 8'hCF},
{8'hFA, 8'hFA, 8'hE8},
{8'hF4, 8'hF5, 8'hEE},
{8'hF6, 8'hF5, 8'hF8},
{8'hF3, 8'hF2, 8'hFD},
{8'hF9, 8'hF8, 8'hFD},
{8'hF7, 8'hF8, 8'hF8},
{8'hED, 8'hEC, 8'hE5},
{8'hE0, 8'hDF, 8'hD3},
{8'hF2, 8'hEF, 8'hE1},
{8'hF8, 8'hF4, 8'hE7},
{8'hF1, 8'hED, 8'hE0},
{8'hF6, 8'hF4, 8'hE8},
{8'hE0, 8'hE0, 8'hD1},
{8'hB9, 8'hBA, 8'hA7},
{8'hD4, 8'hD6, 8'hC1},
{8'h91, 8'h95, 8'h83},
{8'h76, 8'h79, 8'h6F},
{8'h77, 8'h7A, 8'h78},
{8'h76, 8'h7A, 8'h7A},
{8'h93, 8'hA0, 8'h7F},
{8'hD8, 8'hE7, 8'hBD},
{8'hE4, 8'hF1, 8'hCB},
{8'h8A, 8'h92, 8'h84},
{8'h76, 8'h79, 8'h85},
{8'h75, 8'h76, 8'h82},
{8'hB0, 8'hB4, 8'hA3},
{8'hC3, 8'hCB, 8'h9F},
{8'h80, 8'h7F, 8'h7D},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'h7F, 8'h7D, 8'h82},
{8'h7F, 8'h7D, 8'h81},
{8'hFF, 8'hD7, 8'h00},
{8'h7F, 8'h7D, 8'h7F},
{8'h7C, 8'h7A, 8'h7A},
{8'h7F, 8'h7E, 8'h7C},
{8'h95, 8'h94, 8'h91},
{8'h7F, 8'h7F, 8'h7B},
{8'h7C, 8'h7D, 8'h7A},
{8'h84, 8'h82, 8'h78},
{8'h95, 8'h93, 8'h83},
{8'h90, 8'h93, 8'h83},
{8'h7B, 8'h7E, 8'h73},
{8'h7E, 8'h76, 8'h6A},
{8'hB4, 8'h94, 8'h80},
{8'hEF, 8'hC0, 8'hA6},
{8'hED, 8'hCC, 8'hB3},
{8'hEB, 8'hE0, 8'hC3},
{8'hE7, 8'hF1, 8'hD1},
{8'hE2, 8'hF1, 8'hD7},
{8'hF2, 8'hF8, 8'hE4},
{8'hF5, 8'hF4, 8'hE0},
{8'hFA, 8'hF9, 8'hE2},
{8'hF7, 8'hFC, 8'hE3},
{8'hFF, 8'hFB, 8'hFF},
{8'hF6, 8'hF0, 8'hEE},
{8'h76, 8'h7A, 8'h97},
{8'h2B, 8'h50, 8'hAA},
{8'h09, 8'h56, 8'hC8},
{8'h03, 8'h5C, 8'hB4},
{8'h11, 8'h4F, 8'h92},
{8'h13, 8'h24, 8'h70},
{8'h08, 8'h21, 8'h7B},
{8'h18, 8'h49, 8'h9B},
{8'h18, 8'h57, 8'hA4},
{8'h19, 8'h57, 8'hAC},
{8'h1E, 8'h4F, 8'hA9},
{8'h1E, 8'h39, 8'h85},
{8'h01, 8'h06, 8'h2E},
{8'h05, 8'h05, 8'h12},
{8'h00, 8'h09, 8'h1E},
{8'h0B, 8'h00, 8'h01},
{8'h0F, 8'h05, 8'h09},
{8'h1E, 8'h42, 8'h75},
{8'h0F, 8'h59, 8'hBD},
{8'h12, 8'h54, 8'hCC},
{8'h24, 8'h4C, 8'hC8},
{8'h25, 8'h40, 8'hC2},
{8'h35, 8'h39, 8'h87},
{8'h89, 8'h8F, 8'h53},
{8'hDF, 8'hE8, 8'h73},
{8'h69, 8'h78, 8'h68},
{8'h34, 8'h59, 8'hAA},
{8'h1B, 8'h53, 8'h9E},
{8'h44, 8'h73, 8'h9D},
{8'h0B, 8'h1E, 8'h49},
{8'h02, 8'h18, 8'h35},
{8'h09, 8'h23, 8'h45},
{8'h09, 8'h0F, 8'h3F},
{8'h1B, 8'h1A, 8'h54},
{8'h21, 8'h22, 8'h5E},
{8'h00, 8'h0C, 8'h47},
{8'h16, 8'h41, 8'h8E},
{8'h20, 8'h56, 8'hB9},
{8'h27, 8'h53, 8'h9F},
{8'h25, 8'h56, 8'hA1},
{8'h1A, 8'h51, 8'hA4},
{8'h1E, 8'h5D, 8'hB6},
{8'h13, 8'h58, 8'hB5},
{8'h12, 8'h5A, 8'hBA},
{8'h0E, 8'h58, 8'hB9},
{8'h02, 8'h40, 8'h9B},
{8'h52, 8'h56, 8'h56},
{8'hF4, 8'hF7, 8'hE4},
{8'hF6, 8'hFB, 8'hE1},
{8'hEF, 8'hF4, 8'hD5},
{8'hE1, 8'hE9, 8'hCA},
{8'hEF, 8'hF6, 8'hDE},
{8'hF1, 8'hF7, 8'hE9},
{8'hF5, 8'hFC, 8'hF3},
{8'hFA, 8'hFB, 8'hF9},
{8'hFB, 8'hFB, 8'hF8},
{8'hF9, 8'hFA, 8'hF2},
{8'hFA, 8'hFA, 8'hED},
{8'hE8, 8'hE7, 8'hDA},
{8'hD5, 8'hD2, 8'hC6},
{8'hE4, 8'hE0, 8'hD7},
{8'hF2, 8'hED, 8'hE6},
{8'hF5, 8'hF2, 8'hEC},
{8'hFF, 8'hFF, 8'hF5},
{8'hCA, 8'hCB, 8'hBB},
{8'hC8, 8'hCA, 8'hB7},
{8'hD7, 8'hDB, 8'hC9},
{8'h87, 8'h8B, 8'h7C},
{8'h76, 8'h7B, 8'h71},
{8'h9E, 8'hA4, 8'h9B},
{8'hD8, 8'hE7, 8'hBD},
{8'hE6, 8'hF4, 8'hC9},
{8'hC1, 8'hCF, 8'hAA},
{8'h75, 8'h7E, 8'h66},
{8'h79, 8'h80, 8'h72},
{8'hAE, 8'hB2, 8'hA6},
{8'hEB, 8'hF0, 8'hDB},
{8'hA4, 8'hA9, 8'h8F},
{8'h7B, 8'h79, 8'h7A},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'h7F, 8'h7D, 8'h82},
{8'h7F, 8'h7D, 8'h81},
{8'hFF, 8'hD7, 8'h00},
{8'h7F, 8'h7D, 8'h7F},
{8'h7C, 8'h7A, 8'h7A},
{8'h7E, 8'h7D, 8'h7B},
{8'h95, 8'h94, 8'h91},
{8'h8E, 8'h8F, 8'h89},
{8'h99, 8'hA7, 8'h8B},
{8'hDB, 8'hE2, 8'hBF},
{8'hF1, 8'hF2, 8'hCB},
{8'hEF, 8'hF0, 8'hCC},
{8'hDC, 8'hD8, 8'hC0},
{8'hBB, 8'hA6, 8'h92},
{8'hBD, 8'h8D, 8'h77},
{8'hE3, 8'h9B, 8'h80},
{8'hFA, 8'hA3, 8'h92},
{8'hF6, 8'hB5, 8'hA0},
{8'hF7, 8'hD8, 8'hBD},
{8'hFB, 8'hF6, 8'hD8},
{8'hFA, 8'hF5, 8'hDA},
{8'hFD, 8'hF5, 8'hDC},
{8'hFF, 8'hF4, 8'hDA},
{8'hFD, 8'hF6, 8'hDF},
{8'hF9, 8'hF9, 8'hEE},
{8'hFF, 8'hF9, 8'hE6},
{8'hE0, 8'hD6, 8'hD2},
{8'h51, 8'h68, 8'h94},
{8'h17, 8'h5D, 8'hB4},
{8'h07, 8'h5E, 8'hC1},
{8'h1B, 8'h55, 8'hB8},
{8'h2F, 8'h45, 8'hA9},
{8'h12, 8'h3B, 8'h97},
{8'h06, 8'h2F, 8'h85},
{8'h17, 8'h55, 8'hA9},
{8'h17, 8'h53, 8'hAB},
{8'h1D, 8'h4D, 8'hA3},
{8'h1C, 8'h39, 8'h7F},
{8'h03, 8'h08, 8'h2F},
{8'h05, 8'h05, 8'h17},
{8'h00, 8'h0A, 8'h26},
{8'h03, 8'h01, 8'h10},
{8'h05, 8'h02, 8'h1D},
{8'h14, 8'h3B, 8'h7A},
{8'h1C, 8'h5B, 8'hA8},
{8'h2A, 8'h55, 8'h8B},
{8'h56, 8'h69, 8'h81},
{8'h83, 8'h90, 8'h97},
{8'hC8, 8'hBD, 8'h77},
{8'hF0, 8'hD4, 8'h76},
{8'hF0, 8'hBD, 8'h5A},
{8'hEC, 8'hBA, 8'h6B},
{8'hC4, 8'hB1, 8'h83},
{8'h8E, 8'h91, 8'h81},
{8'h55, 8'h5F, 8'h6D},
{8'h1A, 8'h1E, 8'h49},
{8'h1F, 8'h34, 8'hA5},
{8'h21, 8'h3B, 8'hA3},
{8'h01, 8'h11, 8'h4E},
{8'h13, 8'h32, 8'h4B},
{8'h0B, 8'h23, 8'h44},
{8'h0D, 8'h2A, 8'h70},
{8'h21, 8'h4C, 8'h9E},
{8'h0C, 8'h37, 8'h7A},
{8'h10, 8'h22, 8'h56},
{8'h0A, 8'h14, 8'h4D},
{8'h05, 8'h15, 8'h57},
{8'h0A, 8'h2C, 8'h78},
{8'h0F, 8'h43, 8'h95},
{8'h1B, 8'h5A, 8'hB2},
{8'h16, 8'h59, 8'hB5},
{8'h0E, 8'h4C, 8'hA4},
{8'h2A, 8'h29, 8'h43},
{8'hF2, 8'hEB, 8'hF2},
{8'hFA, 8'hF3, 8'hFA},
{8'hFA, 8'hF3, 8'hF2},
{8'hF9, 8'hF3, 8'hEC},
{8'hE8, 8'hDC, 8'hD7},
{8'hEC, 8'hDE, 8'hDC},
{8'hE7, 8'hD9, 8'hDA},
{8'hDF, 8'hE1, 8'hD1},
{8'hEB, 8'hEE, 8'hDB},
{8'hF1, 8'hF3, 8'hDF},
{8'hF2, 8'hF4, 8'hE0},
{8'hEA, 8'hE9, 8'hDB},
{8'hE1, 8'hDE, 8'hD6},
{8'hED, 8'hE7, 8'hE5},
{8'hF7, 8'hF2, 8'hF3},
{8'hE5, 8'hE2, 8'hDB},
{8'hCB, 8'hCA, 8'hBF},
{8'hDD, 8'hDE, 8'hCD},
{8'hD0, 8'hD3, 8'hBC},
{8'hAC, 8'hB2, 8'h96},
{8'h9C, 8'hA2, 8'h85},
{8'hBA, 8'hC2, 8'hA5},
{8'hE6, 8'hF0, 8'hD1},
{8'hDF, 8'hF1, 8'hB7},
{8'hE5, 8'hF5, 8'hC5},
{8'hC3, 8'hD0, 8'hAB},
{8'h82, 8'h8E, 8'h68},
{8'hAF, 8'hBA, 8'h8D},
{8'hEC, 8'hF6, 8'hCC},
{8'hCC, 8'hD1, 8'hBA},
{8'h7C, 8'h7E, 8'h79},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'h7F, 8'h7D, 8'h82},
{8'h7F, 8'h7D, 8'h81},
{8'hFF, 8'hD7, 8'h00},
{8'h7F, 8'h7D, 8'h7F},
{8'h80, 8'h7F, 8'h7E},
{8'h7E, 8'h7D, 8'h7B},
{8'h88, 8'h87, 8'h84},
{8'hAD, 8'hAD, 8'hA6},
{8'hD4, 8'hE3, 8'hB8},
{8'hF3, 8'hFC, 8'hC7},
{8'hE9, 8'hED, 8'hB4},
{8'hEF, 8'hF4, 8'hBE},
{8'hF2, 8'hF7, 8'hCC},
{8'hFC, 8'hF4, 8'hD1},
{8'hF1, 8'hD7, 8'hB2},
{8'hCA, 8'h97, 8'h70},
{8'hEE, 8'h96, 8'h77},
{8'hF8, 8'hA6, 8'h89},
{8'hF9, 8'hAF, 8'h8F},
{8'hFC, 8'hBC, 8'h9E},
{8'hFD, 8'hC2, 8'hA6},
{8'hFB, 8'hC2, 8'hA6},
{8'hF6, 8'hC2, 8'hA5},
{8'hFC, 8'hD7, 8'hB9},
{8'hF6, 8'hFD, 8'hD3},
{8'hFB, 8'hFB, 8'hE4},
{8'hFF, 8'hF3, 8'hDB},
{8'hC1, 8'hB3, 8'h88},
{8'h84, 8'h8C, 8'h7D},
{8'h37, 8'h55, 8'h8E},
{8'h20, 8'h50, 8'hBC},
{8'h19, 8'h52, 8'hC2},
{8'h1B, 8'h55, 8'hAF},
{8'h0F, 8'h46, 8'h9F},
{8'h0B, 8'h44, 8'h9F},
{8'h1B, 8'h54, 8'hAE},
{8'h1E, 8'h4B, 8'h9B},
{8'h10, 8'h28, 8'h64},
{8'h04, 8'h06, 8'h2C},
{8'h05, 8'h05, 8'h1A},
{8'h04, 8'h06, 8'h1E},
{8'h02, 8'h00, 8'h17},
{8'h00, 8'h00, 8'h24},
{8'h24, 8'h44, 8'h68},
{8'h74, 8'h87, 8'h84},
{8'hC3, 8'hB4, 8'h72},
{8'hE9, 8'hD1, 8'h65},
{8'hE1, 8'hD7, 8'h6C},
{8'hE5, 8'hCB, 8'h8E},
{8'hF1, 8'hC7, 8'h79},
{8'hF5, 8'hC7, 8'h97},
{8'hF4, 8'hC2, 8'hBC},
{8'hF1, 8'hCD, 8'h97},
{8'hE7, 8'hDA, 8'h4D},
{8'hDB, 8'hD2, 8'h56},
{8'hA4, 8'h90, 8'h6E},
{8'h6B, 8'h6A, 8'h7F},
{8'h42, 8'h4C, 8'h88},
{8'h1E, 8'h38, 8'h7B},
{8'h0A, 8'h32, 8'h56},
{8'h06, 8'h24, 8'h44},
{8'h13, 8'h33, 8'h70},
{8'h07, 8'h11, 8'h4E},
{8'h02, 8'h03, 8'h24},
{8'h00, 8'h00, 8'h2C},
{8'h05, 8'h0D, 8'h40},
{8'h13, 8'h24, 8'h5D},
{8'h12, 8'h29, 8'h6A},
{8'h0A, 8'h23, 8'h68},
{8'h10, 8'h31, 8'h78},
{8'h16, 8'h42, 8'h8C},
{8'h16, 8'h3E, 8'h84},
{8'h11, 8'h0E, 8'h2A},
{8'hD9, 8'hD2, 8'hE1},
{8'hFF, 8'hFA, 8'hFF},
{8'hFF, 8'hF7, 8'hF3},
{8'hFE, 8'hEF, 8'hE1},
{8'hED, 8'hD7, 8'hC3},
{8'hD9, 8'hBF, 8'hA9},
{8'hCA, 8'hB1, 8'h9A},
{8'hD3, 8'hD5, 8'hBB},
{8'hD0, 8'hD5, 8'hBA},
{8'hE0, 8'hE4, 8'hC9},
{8'hE5, 8'hE7, 8'hD0},
{8'hDE, 8'hDD, 8'hCE},
{8'hF6, 8'hF2, 8'hEC},
{8'hFD, 8'hF9, 8'hFA},
{8'hFD, 8'hF9, 8'hFD},
{8'hC0, 8'hBF, 8'hAE},
{8'hA0, 8'hA0, 8'h8B},
{8'hE5, 8'hE7, 8'hCC},
{8'hE1, 8'hE5, 8'hC3},
{8'hD8, 8'hE0, 8'hB5},
{8'hE7, 8'hEF, 8'hC0},
{8'hE4, 8'hF0, 8'hBA},
{8'hE3, 8'hF1, 8'hB8},
{8'hE3, 8'hF6, 8'hB2},
{8'hE4, 8'hF5, 8'hC0},
{8'hE0, 8'hEE, 8'hC7},
{8'hD8, 8'hE6, 8'hB5},
{8'hE8, 8'hF6, 8'hB6},
{8'hE8, 8'hF5, 8'hBA},
{8'hA1, 8'hA6, 8'h8F},
{8'h78, 8'h78, 8'h81},
{8'h7E, 8'h7C, 8'h80},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'h7F, 8'h7D, 8'h82},
{8'h7F, 8'h7D, 8'h81},
{8'hFF, 8'hD7, 8'h00},
{8'h7F, 8'h7D, 8'h7F},
{8'h7B, 8'h7A, 8'h79},
{8'h83, 8'h82, 8'h80},
{8'h7C, 8'h7B, 8'h78},
{8'hB5, 8'hB5, 8'hAE},
{8'hE7, 8'hF0, 8'hC4},
{8'hF1, 8'hF6, 8'hBE},
{8'hEF, 8'hF4, 8'hB4},
{8'hEC, 8'hF9, 8'hB8},
{8'hE5, 8'hF9, 8'hC3},
{8'hE8, 8'hFA, 8'hC9},
{8'hF2, 8'hF8, 8'hC6},
{8'hEE, 8'hE6, 8'hB0},
{8'hD5, 8'hBC, 8'h80},
{8'hD2, 8'hA3, 8'h6D},
{8'hEB, 8'hA4, 8'h76},
{8'hF3, 8'hA0, 8'h79},
{8'hF2, 8'hA0, 8'h7B},
{8'hEB, 8'hA5, 8'h7E},
{8'hEC, 8'hB3, 8'h8B},
{8'hEC, 8'hBD, 8'h94},
{8'hEF, 8'hDC, 8'hB5},
{8'hFD, 8'hF5, 8'hE1},
{8'hFE, 8'hFB, 8'hE4},
{8'hF9, 8'hE5, 8'hA8},
{8'hFB, 8'hDA, 8'h89},
{8'hCE, 8'hBC, 8'h8B},
{8'h57, 8'h70, 8'h7C},
{8'h19, 8'h5C, 8'h92},
{8'h1B, 8'h57, 8'hAA},
{8'h1A, 8'h54, 8'hAF},
{8'h0F, 8'h48, 8'hA9},
{8'h1C, 8'h4F, 8'hA9},
{8'h26, 8'h4C, 8'h92},
{8'h03, 8'h10, 8'h41},
{8'h01, 8'h03, 8'h23},
{8'h05, 8'h03, 8'h1F},
{8'h07, 8'h00, 8'h31},
{8'h21, 8'h04, 8'h09},
{8'h62, 8'h38, 8'h0C},
{8'hCE, 8'hB6, 8'h64},
{8'hF4, 8'hDA, 8'h78},
{8'hEB, 8'hC7, 8'h63},
{8'hEC, 8'hCE, 8'h88},
{8'hF1, 8'hE7, 8'hC6},
{8'hFC, 8'hFD, 8'hDE},
{8'hFD, 8'hFF, 8'hE6},
{8'hFC, 8'hFE, 8'hEA},
{8'hFA, 8'hFF, 8'hE7},
{8'hFB, 8'hFF, 8'hE7},
{8'hFE, 8'hFD, 8'hE1},
{8'hF5, 8'hED, 8'hC4},
{8'hED, 8'hE0, 8'h9B},
{8'hDA, 8'hDD, 8'h6C},
{8'hB5, 8'hB8, 8'h89},
{8'h77, 8'h7C, 8'h8B},
{8'h1D, 8'h29, 8'h47},
{8'h04, 8'h10, 8'h37},
{8'h07, 8'h0A, 8'h44},
{8'h06, 8'h01, 8'h2F},
{8'h09, 8'h05, 8'h18},
{8'h0F, 8'h30, 8'h73},
{8'h23, 8'h4F, 8'h98},
{8'h28, 8'h58, 8'hA3},
{8'h25, 8'h57, 8'hA5},
{8'h22, 8'h55, 8'hA4},
{8'h20, 8'h50, 8'h9E},
{8'h1D, 8'h4C, 8'h98},
{8'h1D, 8'h49, 8'h90},
{8'h18, 8'h38, 8'h58},
{8'h42, 8'h61, 8'h77},
{8'h92, 8'hAB, 8'hB5},
{8'hBB, 8'hCD, 8'hCB},
{8'hE8, 8'hF0, 8'hE3},
{8'hE6, 8'hEA, 8'hCF},
{8'hE0, 8'hDF, 8'hBC},
{8'hEC, 8'hE8, 8'hC4},
{8'hEA, 8'hEE, 8'hD6},
{8'hE7, 8'hEA, 8'hD2},
{8'hE7, 8'hEB, 8'hD2},
{8'hEB, 8'hEE, 8'hD8},
{8'hFB, 8'hFB, 8'hEC},
{8'hF6, 8'hF3, 8'hEC},
{8'hFA, 8'hF5, 8'hF6},
{8'hFC, 8'hF7, 8'hF9},
{8'hA2, 8'hA2, 8'h88},
{8'hA1, 8'hA3, 8'h84},
{8'hE3, 8'hE7, 8'hC4},
{8'hE8, 8'hED, 8'hC4},
{8'hE8, 8'hF1, 8'hBE},
{8'hE6, 8'hF2, 8'hB4},
{8'hE6, 8'hF5, 8'hB0},
{8'hE2, 8'hF2, 8'hA8},
{8'hE2, 8'hF5, 8'hAE},
{8'hE2, 8'hF4, 8'hBB},
{8'hE3, 8'hF2, 8'hC4},
{8'hE6, 8'hF4, 8'hBF},
{8'hE8, 8'hF6, 8'hB7},
{8'hCE, 8'hD8, 8'hA4},
{8'h7C, 8'h80, 8'h6E},
{8'h7B, 8'h7A, 8'h87},
{8'h7F, 8'h7D, 8'h82},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'h7F, 8'h7D, 8'h82},
{8'h7F, 8'h7D, 8'h81},
{8'hFF, 8'hD7, 8'h00},
{8'h80, 8'h7D, 8'h80},
{8'h82, 8'h80, 8'h80},
{8'h83, 8'h82, 8'h80},
{8'h7C, 8'h7B, 8'h78},
{8'h8C, 8'h8C, 8'h86},
{8'hE0, 8'hE8, 8'hC3},
{8'hF3, 8'hF8, 8'hC6},
{8'hEE, 8'hF2, 8'hB6},
{8'hEF, 8'hFB, 8'hBE},
{8'hE0, 8'hFB, 8'hC1},
{8'hDF, 8'hFD, 8'hC9},
{8'hE7, 8'hFC, 8'hC7},
{8'hE8, 8'hF5, 8'hBC},
{8'hE3, 8'hFB, 8'hB7},
{8'hEF, 8'hEC, 8'hAD},
{8'hD3, 8'hAA, 8'h77},
{8'hE0, 8'h9E, 8'h72},
{8'hF2, 8'hB8, 8'h8C},
{8'hEE, 8'hC6, 8'h99},
{8'hE6, 8'hCA, 8'h9E},
{8'hFC, 8'hEA, 8'hC2},
{8'hF9, 8'hD1, 8'hC1},
{8'hFA, 8'hE4, 8'hD3},
{8'hFC, 8'hFE, 8'hF5},
{8'hFC, 8'hF9, 8'hE6},
{8'hF7, 8'hDC, 8'h94},
{8'hFF, 8'hE8, 8'h6F},
{8'hE0, 8'hDC, 8'h79},
{8'h69, 8'h85, 8'h66},
{8'h1F, 8'h59, 8'hA0},
{8'h1A, 8'h53, 8'hAE},
{8'h14, 8'h48, 8'hAC},
{8'h16, 8'h42, 8'h9B},
{8'h23, 8'h44, 8'h80},
{8'h02, 8'h06, 8'h2B},
{8'h02, 8'h00, 8'h1A},
{8'h08, 8'h01, 8'h1C},
{8'h0C, 8'h00, 8'h10},
{8'h7F, 8'h35, 8'h19},
{8'hE8, 8'h76, 8'h32},
{8'hF3, 8'h9F, 8'h63},
{8'hED, 8'hC7, 8'hA0},
{8'hF9, 8'hEF, 8'hCB},
{8'hFB, 8'hFC, 8'hDB},
{8'hF5, 8'hFF, 8'hEA},
{8'hFB, 8'hFB, 8'hF2},
{8'hF6, 8'hFF, 8'hDB},
{8'hEF, 8'hFF, 8'hD1},
{8'hED, 8'hFF, 8'hE3},
{8'hF4, 8'hFF, 8'hF7},
{8'hFD, 8'hFB, 8'hF7},
{8'hFF, 8'hF8, 8'hF3},
{8'hFF, 8'hF6, 8'hEE},
{8'hF4, 8'hF6, 8'hD4},
{8'hED, 8'hEC, 8'hB7},
{8'hE6, 8'hDB, 8'h9B},
{8'hC1, 8'hA9, 8'h7A},
{8'h3D, 8'h25, 8'h27},
{8'h09, 8'h00, 8'h22},
{8'h07, 8'h06, 8'h22},
{8'h14, 8'h23, 8'h32},
{8'h22, 8'h5D, 8'hAE},
{8'h1B, 8'h5C, 8'hB5},
{8'h10, 8'h54, 8'hB0},
{8'h11, 8'h57, 8'hB6},
{8'h0F, 8'h57, 8'hB5},
{8'h10, 8'h56, 8'hB4},
{8'h14, 8'h57, 8'hB2},
{8'h15, 8'h56, 8'hB0},
{8'h17, 8'h5D, 8'hB4},
{8'h10, 8'h52, 8'hA3},
{8'h0B, 8'h46, 8'h8D},
{8'h14, 8'h44, 8'h7D},
{8'h35, 8'h55, 8'h80},
{8'h60, 8'h79, 8'h97},
{8'hA9, 8'hB9, 8'hC8},
{8'hE3, 8'hF0, 8'hF6},
{8'hFF, 8'hFF, 8'hFE},
{8'hFF, 8'hFF, 8'hFB},
{8'hFD, 8'hFE, 8'hEF},
{8'hF9, 8'hFB, 8'hEA},
{8'hF6, 8'hF6, 8'hE8},
{8'hF3, 8'hF1, 8'hE6},
{8'hF8, 8'hF5, 8'hF0},
{8'hF0, 8'hEC, 8'hE9},
{8'hAE, 8'hAD, 8'h96},
{8'hC6, 8'hC8, 8'hAE},
{8'hDC, 8'hDF, 8'hC3},
{8'hD9, 8'hDD, 8'hBC},
{8'hD8, 8'hE0, 8'hB5},
{8'hDF, 8'hE9, 8'hB4},
{8'hE5, 8'hF2, 8'hB3},
{8'hEA, 8'hFA, 8'hB4},
{8'hE3, 8'hF5, 8'hB4},
{8'hE2, 8'hF4, 8'hB7},
{8'hE3, 8'hF3, 8'hBC},
{8'hE4, 8'hF2, 8'hC0},
{8'hE7, 8'hF1, 8'hC8},
{8'h94, 8'h9B, 8'h7F},
{8'h7A, 8'h7D, 8'h74},
{8'h7D, 8'h7D, 8'h83},
{8'h7E, 8'h7D, 8'h80},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'h7F, 8'h7D, 8'h82},
{8'h7F, 8'h7D, 8'h81},
{8'hFF, 8'hD7, 8'h00},
{8'h7E, 8'h7C, 8'h7E},
{8'h7B, 8'h7A, 8'h79},
{8'h84, 8'h83, 8'h80},
{8'h7C, 8'h7B, 8'h78},
{8'h7B, 8'h7C, 8'h76},
{8'h9D, 8'hAA, 8'h90},
{8'hF1, 8'hFA, 8'hD2},
{8'hF3, 8'hF7, 8'hC2},
{8'hE8, 8'hF2, 8'hB9},
{8'hE9, 8'hFB, 8'hC9},
{8'hE4, 8'hF7, 8'hCA},
{8'hE9, 8'hF2, 8'hC5},
{8'hF6, 8'hF5, 8'hC5},
{8'hEE, 8'hF8, 8'hCB},
{8'hE1, 8'hD2, 8'hAA},
{8'hD3, 8'hA3, 8'h81},
{8'hF1, 8'hC0, 8'h9E},
{8'hFB, 8'hDD, 8'hB8},
{8'hFD, 8'hF4, 8'hD0},
{8'hF0, 8'hDE, 8'hC3},
{8'hF5, 8'hDC, 8'hC9},
{8'hFE, 8'hF2, 8'hD4},
{8'hFD, 8'hF3, 8'hE0},
{8'hF7, 8'hF9, 8'hF3},
{8'hF7, 8'hFB, 8'hF0},
{8'hFD, 8'hF7, 8'hC7},
{8'hF6, 8'hE3, 8'h8A},
{8'hF6, 8'hDE, 8'h7B},
{8'hE5, 8'hD7, 8'h90},
{8'h32, 8'h66, 8'hA3},
{8'h1A, 8'h4F, 8'hAA},
{8'h1B, 8'h48, 8'hAE},
{8'h13, 8'h35, 8'h8E},
{8'h16, 8'h30, 8'h65},
{8'h00, 8'h04, 8'h1E},
{8'h03, 8'h00, 8'h14},
{8'h0B, 8'h00, 8'h17},
{8'h55, 8'h25, 8'h25},
{8'hD0, 8'h81, 8'h5B},
{8'hF5, 8'hAC, 8'h6E},
{8'hFB, 8'hE9, 8'hB9},
{8'hF9, 8'hFE, 8'hE1},
{8'hFD, 8'hFF, 8'hE2},
{8'hF7, 8'hFB, 8'hE1},
{8'hF7, 8'hFD, 8'hF4},
{8'hFF, 8'hF6, 8'hF3},
{8'hFF, 8'hFA, 8'hE9},
{8'hFC, 8'hFF, 8'hDE},
{8'hFA, 8'hFE, 8'hD7},
{8'hF8, 8'hF7, 8'hD5},
{8'hFF, 8'hFC, 8'hDE},
{8'hFF, 8'hFE, 8'hD7},
{8'hFA, 8'hFD, 8'hCD},
{8'hF8, 8'hFA, 8'hEA},
{8'hFE, 8'hFC, 8'hE9},
{8'hFC, 8'hF5, 8'hE1},
{8'hFC, 8'hEA, 8'hCE},
{8'h9E, 8'h91, 8'h67},
{8'h0D, 8'h12, 8'h01},
{8'h00, 8'h01, 8'h0C},
{8'h19, 8'h29, 8'h79},
{8'h22, 8'h3F, 8'h82},
{8'h0F, 8'h2F, 8'h71},
{8'h03, 8'h21, 8'h6A},
{8'h09, 8'h30, 8'h80},
{8'h18, 8'h54, 8'hAB},
{8'h16, 8'h58, 8'hB3},
{8'h14, 8'h58, 8'hB5},
{8'h13, 8'h59, 8'hB8},
{8'h14, 8'h5C, 8'hC9},
{8'h18, 8'h5A, 8'hC5},
{8'h1D, 8'h55, 8'hB7},
{8'h21, 8'h4B, 8'hA0},
{8'h1A, 8'h34, 8'h7A},
{8'h16, 8'h23, 8'h59},
{8'h09, 8'h0D, 8'h36},
{8'h29, 8'h2A, 8'h48},
{8'h60, 8'h5E, 8'h63},
{8'hAA, 8'hA8, 8'hA6},
{8'hD1, 8'hD0, 8'hC8},
{8'hF7, 8'hF5, 8'hE7},
{8'hF7, 8'hF5, 8'hE4},
{8'hFD, 8'hF9, 8'hE8},
{8'hFF, 8'hFC, 8'hEE},
{8'hCA, 8'hC5, 8'hB8},
{8'hD3, 8'hCF, 8'hC4},
{8'hFB, 8'hF9, 8'hEF},
{8'hFE, 8'hFD, 8'hF2},
{8'hF8, 8'hF8, 8'hEB},
{8'hF2, 8'hF5, 8'hE2},
{8'hD7, 8'hDC, 8'hBE},
{8'hCD, 8'hD7, 8'hAD},
{8'hDF, 8'hEC, 8'hBA},
{8'hE3, 8'hF4, 8'hBC},
{8'hE2, 8'hF5, 8'hB4},
{8'hE3, 8'hF5, 8'hB5},
{8'hE6, 8'hF4, 8'hC8},
{8'hC3, 8'hCB, 8'hBC},
{8'h76, 8'h79, 8'h7C},
{8'h85, 8'h86, 8'h87},
{8'h7E, 8'h80, 8'h77},
{8'h7E, 8'h7D, 8'h7F},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'h7F, 8'h7D, 8'h81},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'h7F, 8'h7E, 8'h7F},
{8'h7F, 8'h7D, 8'h7F},
{8'h7F, 8'h7D, 8'h7F},
{8'h7E, 8'h7C, 8'h7F},
{8'h7C, 8'h7B, 8'h7C},
{8'h7C, 8'h7A, 8'h7A},
{8'h84, 8'h82, 8'h81},
{8'h7C, 8'h7C, 8'h79},
{8'hB5, 8'hC3, 8'hB0},
{8'hB7, 8'hC0, 8'hA2},
{8'hE2, 8'hE7, 8'hBF},
{8'hE0, 8'hE6, 8'hB8},
{8'hB8, 8'hC1, 8'h96},
{8'hC7, 8'hCE, 8'hA6},
{8'hEE, 8'hEE, 8'hC3},
{8'hF8, 8'hEE, 8'hC2},
{8'hFA, 8'hE4, 8'hCB},
{8'hE3, 8'hC1, 8'hAC},
{8'hF9, 8'hD1, 8'hBF},
{8'hF9, 8'hE8, 8'hD3},
{8'hFD, 8'hF9, 8'hE2},
{8'hFF, 8'hF8, 8'hE2},
{8'hFF, 8'hF2, 8'hE4},
{8'hF2, 8'hD0, 8'hC2},
{8'hEA, 8'hCF, 8'h95},
{8'hFB, 8'hE3, 8'hC5},
{8'hFE, 8'hF3, 8'hE6},
{8'hF8, 8'hF8, 8'hE0},
{8'hF6, 8'hFE, 8'hDE},
{8'hF9, 8'hF8, 8'hD8},
{8'hF7, 8'hDA, 8'hA6},
{8'hEF, 8'hCE, 8'h8A},
{8'h2F, 8'h64, 8'hA6},
{8'h1D, 8'h4F, 8'hAB},
{8'h26, 8'h47, 8'hA0},
{8'h0E, 8'h1F, 8'h61},
{8'h03, 8'h0A, 8'h33},
{8'h01, 8'h03, 8'h1E},
{8'h06, 8'h01, 8'h13},
{8'h3A, 8'h22, 8'h2D},
{8'hDD, 8'h9B, 8'h65},
{8'hF9, 8'hC5, 8'h8B},
{8'hFB, 8'hF2, 8'hC7},
{8'hEA, 8'hFF, 8'hEF},
{8'hE7, 8'hFE, 8'hE8},
{8'hFC, 8'hFE, 8'hDB},
{8'hFE, 8'hF8, 8'hDC},
{8'hF8, 8'hF1, 8'hE9},
{8'hF8, 8'hF2, 8'hE1},
{8'hF8, 8'hF4, 8'hDD},
{8'hF9, 8'hF6, 8'hD8},
{8'hF8, 8'hF5, 8'hD5},
{8'hF2, 8'hEA, 8'hDA},
{8'hEE, 8'hE7, 8'hDE},
{8'hF9, 8'hFD, 8'hE2},
{8'hF1, 8'hFF, 8'hCE},
{8'hFD, 8'hFA, 8'hEC},
{8'hFE, 8'hFE, 8'hD3},
{8'hFA, 8'hFD, 8'hCA},
{8'hF2, 8'hF5, 8'hE5},
{8'hE8, 8'hEC, 8'hF6},
{8'h9F, 8'hA7, 8'hB4},
{8'h34, 8'h3A, 8'h51},
{8'h07, 8'h11, 8'h3A},
{8'h04, 8'h01, 8'h26},
{8'h00, 8'h00, 8'h2D},
{8'h0A, 8'h18, 8'h59},
{8'h22, 8'h43, 8'h8F},
{8'h25, 8'h52, 8'hA0},
{8'h23, 8'h56, 8'hA4},
{8'h21, 8'h55, 8'hA6},
{8'h22, 8'h54, 8'hA7},
{8'h1F, 8'h47, 8'h8C},
{8'h12, 8'h35, 8'h74},
{8'h07, 8'h1D, 8'h53},
{8'h03, 8'h0C, 8'h39},
{8'h00, 8'h04, 8'h28},
{8'h02, 8'h05, 8'h23},
{8'h09, 8'h0A, 8'h24},
{8'h0E, 8'h0C, 8'h27},
{8'h00, 8'h0B, 8'h2F},
{8'h00, 8'h0F, 8'h2F},
{8'h12, 8'h24, 8'h40},
{8'h34, 8'h45, 8'h5D},
{8'h66, 8'h73, 8'h84},
{8'h9A, 8'hA3, 8'hB1},
{8'hB0, 8'hB6, 8'hC3},
{8'hB7, 8'hBD, 8'hC9},
{8'hD3, 8'hE0, 8'hE6},
{8'hDD, 8'hE8, 8'hEF},
{8'hE9, 8'hF2, 8'hF9},
{8'hF4, 8'hFA, 8'hFC},
{8'hFF, 8'hFF, 8'hFD},
{8'hFB, 8'hFE, 8'hE8},
{8'hE7, 8'hEC, 8'hC7},
{8'hD3, 8'hDA, 8'hAB},
{8'hDE, 8'hED, 8'hB4},
{8'hE6, 8'hF6, 8'hB4},
{8'hE7, 8'hF3, 8'hB3},
{8'hE6, 8'hEC, 8'hC5},
{8'h92, 8'h93, 8'h8F},
{8'h7D, 8'h7A, 8'h89},
{8'h7E, 8'h7C, 8'h87},
{8'h7B, 8'h7C, 8'h7B},
{8'h82, 8'h7C, 8'h7E},
{8'h81, 8'h7C, 8'h7D},
{8'h80, 8'h7D, 8'h7F},
{8'h80, 8'h7E, 8'h82},
{8'h7F, 8'h7D, 8'h84},
{8'h80, 8'h7C, 8'h82},
{8'h81, 8'h7C, 8'h7E},
{8'h82, 8'h7D, 8'h7A},
{8'h7E, 8'h7E, 8'h7E},
{8'h7E, 8'h7E, 8'h7E},
{8'h7F, 8'h7E, 8'h7E},
{8'h7F, 8'h7E, 8'h7E},
{8'h7F, 8'h7E, 8'h7E},
{8'h7E, 8'h7E, 8'h7F},
{8'h7E, 8'h7E, 8'h7F},
{8'h7D, 8'h7E, 8'h80},
{8'h7F, 8'h7D, 8'h7F},
{8'h7F, 8'h7D, 8'h7F},
{8'h7F, 8'h7D, 8'h7F},
{8'h80, 8'h7D, 8'h7F},
{8'h80, 8'h7C, 8'h7F},
{8'h80, 8'h7C, 8'h7F},
{8'h81, 8'h7C, 8'h7F},
{8'h81, 8'h7C, 8'h7F},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'h7F, 8'h7F, 8'h77},
{8'h7F, 8'h7E, 8'h79},
{8'h7F, 8'h7D, 8'h7E},
{8'h7E, 8'h7C, 8'h81},
{8'h7E, 8'h7B, 8'h82},
{8'h7E, 8'h7C, 8'h81},
{8'h81, 8'h7E, 8'h81},
{8'h93, 8'h92, 8'h90},
{8'hCE, 8'hCE, 8'hBE},
{8'h78, 8'h7A, 8'h67},
{8'h85, 8'h89, 8'h73},
{8'hD8, 8'hDD, 8'hC0},
{8'hED, 8'hF5, 8'hD0},
{8'hEB, 8'hF4, 8'hC6},
{8'hEC, 8'hF8, 8'hC1},
{8'hF0, 8'hFC, 8'hC2},
{8'hE9, 8'hD0, 8'hAE},
{8'hE4, 8'hD9, 8'hBC},
{8'hF3, 8'hFC, 8'hE4},
{8'hF0, 8'hFF, 8'hED},
{8'hF6, 8'hFD, 8'hEE},
{8'hFB, 8'hF7, 8'hE5},
{8'hFF, 8'hFA, 8'hE1},
{8'hFB, 8'hF0, 8'hCE},
{8'hFA, 8'hBD, 8'h87},
{8'hF5, 8'hB2, 8'h84},
{8'hFE, 8'hD8, 8'hB8},
{8'hFD, 8'hF7, 8'hE5},
{8'hEF, 8'hFF, 8'hF2},
{8'hF2, 8'hFF, 8'hE8},
{8'hFD, 8'hED, 8'hBE},
{8'hC5, 8'h9C, 8'h6A},
{8'h18, 8'h55, 8'hAD},
{8'h24, 8'h4E, 8'hAD},
{8'h30, 8'h3B, 8'h70},
{8'h04, 8'h04, 8'h0D},
{8'h00, 8'h01, 8'h11},
{8'h01, 8'h01, 8'h2C},
{8'h04, 8'h00, 8'h11},
{8'h6E, 8'h54, 8'h3D},
{8'hFF, 8'hC2, 8'h8B},
{8'hFA, 8'hE2, 8'hBC},
{8'hFD, 8'hFF, 8'hEB},
{8'hF4, 8'hFA, 8'hE9},
{8'hF9, 8'hF6, 8'hDD},
{8'hF9, 8'hF0, 8'hD8},
{8'hF8, 8'hF1, 8'hE8},
{8'hF7, 8'hF6, 8'hF8},
{8'hF8, 8'hF6, 8'hF8},
{8'hF8, 8'hF6, 8'hF5},
{8'hF9, 8'hF6, 8'hF1},
{8'hF9, 8'hF5, 8'hEB},
{8'hF4, 8'hF0, 8'hE0},
{8'hF2, 8'hEB, 8'hD5},
{8'hEE, 8'hE5, 8'hCC},
{8'hFF, 8'hFA, 8'hDF},
{8'hFF, 8'hFC, 8'hE5},
{8'hFA, 8'hF9, 8'hE6},
{8'hED, 8'hEE, 8'hDE},
{8'hED, 8'hF2, 8'hE5},
{8'hF6, 8'hFB, 8'hF6},
{8'hFF, 8'hFF, 8'hFF},
{8'hF4, 8'hF3, 8'hF5},
{8'h92, 8'h91, 8'h96},
{8'h15, 8'h22, 8'h3C},
{8'h19, 8'h30, 8'h6E},
{8'h28, 8'h50, 8'hB4},
{8'h1C, 8'h54, 8'hC0},
{8'h18, 8'h57, 8'hB1},
{8'h17, 8'h50, 8'h98},
{8'h18, 8'h3C, 8'h85},
{8'h10, 8'h27, 8'h74},
{8'h0D, 8'h23, 8'h50},
{8'h08, 8'h23, 8'h55},
{8'h0E, 8'h2E, 8'h6B},
{8'h16, 8'h3A, 8'h82},
{8'h16, 8'h41, 8'h90},
{8'h12, 8'h46, 8'h98},
{8'h13, 8'h4D, 8'h9E},
{8'h14, 8'h52, 8'hA2},
{8'h0F, 8'h53, 8'hB0},
{8'h0F, 8'h55, 8'hB7},
{8'h0F, 8'h55, 8'hB9},
{8'h0F, 8'h51, 8'hB6},
{8'h11, 8'h4D, 8'hB2},
{8'h0D, 8'h3F, 8'hA2},
{8'h12, 8'h3D, 8'h9E},
{8'h21, 8'h48, 8'hA4},
{8'h1F, 8'h54, 8'h95},
{8'h24, 8'h55, 8'h96},
{8'h30, 8'h58, 8'h99},
{8'h3C, 8'h58, 8'h92},
{8'h52, 8'h6B, 8'h97},
{8'h86, 8'h9C, 8'hB2},
{8'h9E, 8'hB0, 8'hB2},
{8'hBE, 8'hCF, 8'hC1},
{8'hC4, 8'hDD, 8'h97},
{8'hE5, 8'hF7, 8'hB4},
{8'hF1, 8'hFA, 8'hC1},
{8'hCB, 8'hCD, 8'hA3},
{8'h7F, 8'h7C, 8'h66},
{8'h82, 8'h7E, 8'h7D},
{8'h7F, 8'h7C, 8'h90},
{8'h77, 8'h75, 8'h93},
{8'h83, 8'h75, 8'h8F},
{8'h85, 8'h7C, 8'h88},
{8'h80, 8'h80, 8'h7D},
{8'h7A, 8'h7F, 8'h79},
{8'h7A, 8'h7F, 8'h81},
{8'h7E, 8'h7D, 8'h84},
{8'h82, 8'h7C, 8'h7D},
{8'h84, 8'h7D, 8'h76},
{8'h7D, 8'h7F, 8'h7C},
{8'h7D, 8'h7F, 8'h7C},
{8'h7E, 8'h7F, 8'h7A},
{8'h7F, 8'h7E, 8'h7A},
{8'h7F, 8'h7E, 8'h7A},
{8'h7E, 8'h7F, 8'h7B},
{8'h7C, 8'h7F, 8'h7E},
{8'h7B, 8'h7F, 8'h80},
{8'h7E, 8'h7E, 8'h7F},
{8'h7F, 8'h7D, 8'h7F},
{8'h7F, 8'h7D, 8'h7F},
{8'h81, 8'h7C, 8'h7F},
{8'h82, 8'h7C, 8'h7F},
{8'h83, 8'h7C, 8'h7F},
{8'h84, 8'h7B, 8'h7F},
{8'h84, 8'h7B, 8'h7F},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'h7F, 8'h7E, 8'h7C},
{8'h7F, 8'h7E, 8'h7D},
{8'h7F, 8'h7D, 8'h81},
{8'h7F, 8'h7C, 8'h82},
{8'h81, 8'h7F, 8'h84},
{8'h80, 8'h7E, 8'h80},
{8'h78, 8'h77, 8'h74},
{8'hAF, 8'hAE, 8'hA7},
{8'hD3, 8'hD5, 8'hBC},
{8'h80, 8'h84, 8'h66},
{8'hB7, 8'hBB, 8'h9D},
{8'hEA, 8'hEF, 8'hCC},
{8'hF0, 8'hF7, 8'hCF},
{8'hE9, 8'hF1, 8'hC4},
{8'hED, 8'hF7, 8'hC5},
{8'hE5, 8'hEC, 8'hBA},
{8'hE1, 8'hD0, 8'hB3},
{8'hF6, 8'hEE, 8'hD3},
{8'hF0, 8'hEF, 8'hD3},
{8'hFA, 8'hFA, 8'hE1},
{8'hFC, 8'hFA, 8'hE4},
{8'hFB, 8'hF3, 8'hDE},
{8'hFC, 8'hF6, 8'hDF},
{8'hFF, 8'hFC, 8'hE3},
{8'hFB, 8'hE6, 8'hC7},
{8'hEB, 8'hC3, 8'hA3},
{8'hEC, 8'hC2, 8'hA2},
{8'hFE, 8'hEF, 8'hCF},
{8'hFD, 8'hFC, 8'hE1},
{8'hF9, 8'hFD, 8'hE5},
{8'hFE, 8'hFA, 8'hE7},
{8'h86, 8'h78, 8'h6E},
{8'h15, 8'h4D, 8'h9D},
{8'h0B, 8'h27, 8'h79},
{8'h07, 8'h0B, 8'h39},
{8'h06, 8'h08, 8'h15},
{8'h02, 8'h04, 8'h18},
{8'h04, 8'h01, 8'h2C},
{8'h00, 8'h00, 8'h0F},
{8'h6B, 8'h54, 8'h44},
{8'hFD, 8'hCD, 8'hA4},
{8'hFF, 8'hF1, 8'hD5},
{8'hFB, 8'hF7, 8'hE8},
{8'hEF, 8'hF4, 8'hE5},
{8'hF6, 8'hF6, 8'hE3},
{8'hFE, 8'hFB, 8'hE8},
{8'hFE, 8'hFD, 8'hF6},
{8'hFD, 8'hFF, 8'hFF},
{8'hFF, 8'hFF, 8'hFE},
{8'hFF, 8'hFF, 8'hFD},
{8'hFF, 8'hFF, 8'hFA},
{8'hFF, 8'hFF, 8'hF7},
{8'hFD, 8'hFD, 8'hF1},
{8'hFC, 8'hFB, 8'hEB},
{8'hE8, 8'hE3, 8'hD1},
{8'hE4, 8'hE1, 8'hCE},
{8'hF4, 8'hF0, 8'hE0},
{8'hF1, 8'hEE, 8'hDF},
{8'hF8, 8'hFA, 8'hED},
{8'hFD, 8'hFF, 8'hF7},
{8'hFA, 8'hFE, 8'hF8},
{8'hF6, 8'hFA, 8'hF6},
{8'hFE, 8'hFF, 8'hFF},
{8'hFF, 8'hFF, 8'hFF},
{8'hC0, 8'hCF, 8'hD8},
{8'h43, 8'h61, 8'h8A},
{8'h1D, 8'h4B, 8'h99},
{8'h11, 8'h50, 8'hAC},
{8'h08, 8'h4E, 8'hA3},
{8'h07, 8'h45, 8'h92},
{8'h0E, 8'h43, 8'h94},
{8'h18, 8'h4B, 8'hA4},
{8'h10, 8'h51, 8'hBC},
{8'h18, 8'h5B, 8'hC5},
{8'h1B, 8'h5D, 8'hC5},
{8'h16, 8'h57, 8'hBE},
{8'h15, 8'h56, 8'hBD},
{8'h15, 8'h55, 8'hBC},
{8'h15, 8'h53, 8'hBC},
{8'h15, 8'h53, 8'hBA},
{8'h1C, 8'h57, 8'hA7},
{8'h1A, 8'h57, 8'hA7},
{8'h17, 8'h59, 8'hAD},
{8'h16, 8'h5A, 8'hB3},
{8'h13, 8'h58, 8'hB4},
{8'h18, 8'h5A, 8'hB7},
{8'h1A, 8'h5A, 8'hB5},
{8'h19, 8'h56, 8'hB1},
{8'h1B, 8'h55, 8'hB4},
{8'h19, 8'h52, 8'hB7},
{8'h16, 8'h4F, 8'hB8},
{8'h14, 8'h4D, 8'hB7},
{8'h10, 8'h4A, 8'hAF},
{8'h12, 8'h4E, 8'hA7},
{8'h0F, 8'h4E, 8'h9B},
{8'h1B, 8'h59, 8'h9B},
{8'h38, 8'h5E, 8'h77},
{8'h70, 8'h8E, 8'hA0},
{8'hB2, 8'hC8, 8'hD1},
{8'h88, 8'h96, 8'h97},
{8'h7B, 8'h82, 8'h7E},
{8'h7D, 8'h81, 8'h79},
{8'h7F, 8'h83, 8'h79},
{8'h7B, 8'h80, 8'h79},
{8'h77, 8'h7B, 8'h8F},
{8'h78, 8'h7F, 8'h85},
{8'h79, 8'h84, 8'h78},
{8'h7A, 8'h85, 8'h77},
{8'h77, 8'h81, 8'h7F},
{8'h77, 8'h80, 8'h88},
{8'h77, 8'h7F, 8'h8A},
{8'h78, 8'h80, 8'h87},
{8'h7F, 8'h7D, 8'h83},
{8'h81, 8'h7C, 8'h81},
{8'h82, 8'h7C, 8'h80},
{8'h82, 8'h7C, 8'h7F},
{8'h83, 8'h7C, 8'h7E},
{8'h83, 8'h7C, 8'h7E},
{8'h82, 8'h7C, 8'h7F},
{8'h82, 8'h7C, 8'h7F},
{8'h7E, 8'h7E, 8'h80},
{8'h7E, 8'h7E, 8'h80},
{8'h7E, 8'h7E, 8'h80},
{8'h7E, 8'h7E, 8'h80},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'h7F, 8'h7D, 8'h82},
{8'h7F, 8'h7D, 8'h82},
{8'h7F, 8'h7C, 8'h83},
{8'h7F, 8'h7B, 8'h83},
{8'h80, 8'h7E, 8'h82},
{8'h83, 8'h81, 8'h7F},
{8'h81, 8'h80, 8'h78},
{8'hD5, 8'hD7, 8'hC8},
{8'hF0, 8'hF6, 8'hD0},
{8'hD6, 8'hDD, 8'hB3},
{8'hED, 8'hF3, 8'hCA},
{8'hED, 8'hF2, 8'hC8},
{8'hEF, 8'hF6, 8'hCA},
{8'hED, 8'hF3, 8'hC7},
{8'hF0, 8'hF6, 8'hCB},
{8'hD9, 8'hDD, 8'hB6},
{8'hEE, 8'hEA, 8'hD4},
{8'hFF, 8'hFA, 8'hE2},
{8'hFD, 8'hEF, 8'hD4},
{8'hF8, 8'hE5, 8'hC8},
{8'hFF, 8'hF9, 8'hDD},
{8'hFF, 8'hF9, 8'hE0},
{8'hFB, 8'hF4, 8'hE0},
{8'hFA, 8'hF9, 8'hE9},
{8'hFA, 8'hFE, 8'hF1},
{8'hF4, 8'hE8, 8'hD6},
{8'hF0, 8'hD1, 8'hB7},
{8'hFC, 8'hE6, 8'hC4},
{8'hFF, 8'hF8, 8'hD8},
{8'hFF, 8'hFA, 8'hEA},
{8'hEF, 8'hF1, 8'hF6},
{8'h68, 8'h70, 8'h8A},
{8'h2C, 8'h56, 8'h9A},
{8'h1A, 8'h36, 8'h76},
{8'h00, 8'h03, 8'h2A},
{8'h06, 8'h06, 8'h19},
{8'h02, 8'h02, 8'h1C},
{8'h07, 8'h02, 8'h2A},
{8'h01, 8'h00, 8'h11},
{8'h54, 8'h44, 8'h3C},
{8'hF0, 8'hC9, 8'hB2},
{8'hFC, 8'hE1, 8'hD3},
{8'hF9, 8'hF0, 8'hE7},
{8'hFD, 8'hFF, 8'hF7},
{8'hFD, 8'hFE, 8'hF3},
{8'hFE, 8'hFE, 8'hF4},
{8'hFD, 8'hFD, 8'hFA},
{8'hF9, 8'hFF, 8'hFF},
{8'hFB, 8'hFF, 8'hFB},
{8'hFD, 8'hFF, 8'hFA},
{8'hFD, 8'hFE, 8'hFA},
{8'hFD, 8'hFE, 8'hF9},
{8'hFA, 8'hFA, 8'hF5},
{8'hFC, 8'hFC, 8'hF6},
{8'hFD, 8'hFD, 8'hF8},
{8'hDF, 8'hDE, 8'hD7},
{8'hD2, 8'hCA, 8'hC4},
{8'hFA, 8'hF7, 8'hF0},
{8'hFD, 8'hFE, 8'hF7},
{8'hFC, 8'hFE, 8'hF8},
{8'hFB, 8'hFE, 8'hF9},
{8'hF9, 8'hFC, 8'hF6},
{8'hF9, 8'hFB, 8'hF5},
{8'hFC, 8'hFC, 8'hF7},
{8'hFA, 8'hFF, 8'hFD},
{8'hD2, 8'hE6, 8'hEB},
{8'h43, 8'h6B, 8'h9A},
{8'h0F, 8'h4C, 8'h95},
{8'h0F, 8'h57, 8'hA6},
{8'h12, 8'h5D, 8'hAF},
{8'h16, 8'h5B, 8'hB3},
{8'h18, 8'h57, 8'hB6},
{8'h10, 8'h57, 8'hC5},
{8'h11, 8'h58, 8'hC3},
{8'h14, 8'h58, 8'hBD},
{8'h17, 8'h59, 8'hB7},
{8'h1A, 8'h58, 8'hB2},
{8'h1B, 8'h57, 8'hAF},
{8'h1C, 8'h53, 8'hAB},
{8'h1C, 8'h51, 8'hA9},
{8'h1F, 8'h57, 8'hA3},
{8'h14, 8'h4E, 8'h9D},
{8'h0E, 8'h4F, 8'hA2},
{8'h12, 8'h5A, 8'hB1},
{8'h0F, 8'h5B, 8'hB5},
{8'h0A, 8'h57, 8'hB1},
{8'h0A, 8'h57, 8'hB1},
{8'h0F, 8'h5B, 8'hB4},
{8'h14, 8'h57, 8'hBA},
{8'h14, 8'h56, 8'hBD},
{8'h16, 8'h55, 8'hBC},
{8'h1A, 8'h53, 8'hBB},
{8'h1B, 8'h50, 8'hB2},
{8'h16, 8'h46, 8'h9E},
{8'h0E, 8'h3B, 8'h86},
{8'h04, 8'h2E, 8'h75},
{8'h0C, 8'h1D, 8'h7E},
{8'h0F, 8'h1B, 8'h76},
{8'h1F, 8'h27, 8'h6F},
{8'h2E, 8'h32, 8'h64},
{8'h53, 8'h53, 8'h6E},
{8'h74, 8'h72, 8'h7A},
{8'h81, 8'h7E, 8'h78},
{8'h86, 8'h84, 8'h74},
{8'h7F, 8'h8A, 8'h69},
{8'h7F, 8'h88, 8'h69},
{8'h80, 8'h81, 8'h70},
{8'h81, 8'h7B, 8'h80},
{8'h83, 8'h78, 8'h91},
{8'h81, 8'h79, 8'h92},
{8'h7C, 8'h7E, 8'h84},
{8'h7B, 8'h81, 8'h77},
{8'h80, 8'h7C, 8'h83},
{8'h81, 8'h7B, 8'h84},
{8'h81, 8'h7B, 8'h84},
{8'h82, 8'h7B, 8'h83},
{8'h83, 8'h7B, 8'h83},
{8'h85, 8'h7B, 8'h81},
{8'h86, 8'h7A, 8'h7F},
{8'h86, 8'h7A, 8'h7E},
{8'h80, 8'h7D, 8'h80},
{8'h7E, 8'h7D, 8'h80},
{8'h7E, 8'h7E, 8'h80},
{8'h7D, 8'h7E, 8'h80},
{8'h7C, 8'h7E, 8'h80},
{8'h7B, 8'h7F, 8'h80},
{8'h7B, 8'h80, 8'h80},
{8'h7A, 8'h80, 8'h80},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'h7F, 8'h7C, 8'h83},
{8'h7F, 8'h7C, 8'h85},
{8'h7F, 8'h7C, 8'h85},
{8'h80, 8'h7D, 8'h85},
{8'h83, 8'h81, 8'h84},
{8'h7C, 8'h7B, 8'h78},
{8'h79, 8'h79, 8'h6E},
{8'hC4, 8'hC6, 8'hB4},
{8'hF1, 8'hF8, 8'hCB},
{8'hEF, 8'hF6, 8'hC5},
{8'hEF, 8'hF7, 8'hC4},
{8'hE5, 8'hEB, 8'hBA},
{8'hD7, 8'hDB, 8'hAC},
{8'hD9, 8'hDB, 8'hB2},
{8'hCE, 8'hCF, 8'hAC},
{8'hDB, 8'hDD, 8'hBE},
{8'hFA, 8'hFD, 8'hE9},
{8'hFE, 8'hF6, 8'hE0},
{8'hFE, 8'hE2, 8'hCA},
{8'hEA, 8'hBC, 8'h9F},
{8'hFB, 8'hDF, 8'hC0},
{8'hFF, 8'hF6, 8'hDA},
{8'hFF, 8'hFA, 8'hE8},
{8'hFE, 8'hFD, 8'hF0},
{8'hF4, 8'hF9, 8'hE7},
{8'hFA, 8'hF9, 8'hE9},
{8'hFF, 8'hFA, 8'hEA},
{8'hFD, 8'hF2, 8'hDE},
{8'hFE, 8'hF5, 8'hE0},
{8'hFF, 8'hF8, 8'hF0},
{8'hE1, 8'hDE, 8'hEE},
{8'h55, 8'h59, 8'h7F},
{8'h1A, 8'h2E, 8'h5F},
{8'h04, 8'h11, 8'h39},
{8'h01, 8'h03, 8'h1E},
{8'h03, 8'h06, 8'h1F},
{8'h04, 8'h00, 8'h21},
{8'h06, 8'h01, 8'h23},
{8'h05, 8'h01, 8'h15},
{8'h2E, 8'h27, 8'h2C},
{8'hC6, 8'hA3, 8'hA1},
{8'hF6, 8'hDF, 8'hDD},
{8'hFF, 8'hFC, 8'hFA},
{8'hFF, 8'hFA, 8'hF8},
{8'hFF, 8'hFF, 8'hFC},
{8'hFD, 8'hFE, 8'hFD},
{8'hFB, 8'hFE, 8'hFF},
{8'hFA, 8'hFE, 8'hFF},
{8'hFD, 8'hFF, 8'hFA},
{8'hFD, 8'hFE, 8'hFA},
{8'hFD, 8'hFE, 8'hFB},
{8'hFD, 8'hFE, 8'hFC},
{8'hFE, 8'hFE, 8'hFE},
{8'hFC, 8'hFB, 8'hFC},
{8'hFB, 8'hFB, 8'hFC},
{8'hFA, 8'hF9, 8'hFA},
{8'hD0, 8'hC4, 8'hC7},
{8'hE9, 8'hE0, 8'hE1},
{8'hFF, 8'hFF, 8'hFD},
{8'hFD, 8'hFD, 8'hF8},
{8'hFC, 8'hFE, 8'hF8},
{8'hFD, 8'hFD, 8'hF7},
{8'hFE, 8'hFE, 8'hF7},
{8'hFE, 8'hFC, 8'hF4},
{8'hFE, 8'hFA, 8'hF0},
{8'hFF, 8'hFF, 8'hFF},
{8'hD0, 8'hE5, 8'hEF},
{8'h3D, 8'h66, 8'h9A},
{8'h1C, 8'h52, 8'h98},
{8'h1A, 8'h54, 8'hA5},
{8'h1B, 8'h54, 8'hAB},
{8'h1A, 8'h50, 8'hA8},
{8'h25, 8'h51, 8'h92},
{8'h20, 8'h4B, 8'h8E},
{8'h17, 8'h43, 8'h8B},
{8'h0E, 8'h35, 8'h81},
{8'h0B, 8'h30, 8'h7B},
{8'h05, 8'h2C, 8'h70},
{8'h05, 8'h2A, 8'h67},
{8'h0D, 8'h2C, 8'h66},
{8'h08, 8'h35, 8'h8D},
{8'h07, 8'h45, 8'hA1},
{8'h11, 8'h56, 8'hB4},
{8'h0E, 8'h57, 8'hB5},
{8'h0F, 8'h57, 8'hB5},
{8'h12, 8'h5A, 8'hB4},
{8'h15, 8'h5B, 8'hB1},
{8'h16, 8'h5B, 8'hAE},
{8'h1A, 8'h5B, 8'hA8},
{8'h15, 8'h4F, 8'h9B},
{8'h12, 8'h3D, 8'h87},
{8'h13, 8'h30, 8'h71},
{8'h07, 8'h18, 8'h50},
{8'h03, 8'h08, 8'h32},
{8'h01, 8'h00, 8'h1C},
{8'h04, 8'h00, 8'h13},
{8'h00, 8'h06, 8'h0D},
{8'h00, 8'h05, 8'h0E},
{8'h00, 8'h03, 8'h10},
{8'h00, 8'h02, 8'h17},
{8'h00, 8'h00, 8'h1B},
{8'h14, 8'h15, 8'h39},
{8'h3C, 8'h41, 8'h6C},
{8'h51, 8'h55, 8'h84},
{8'h4C, 8'h50, 8'h76},
{8'h63, 8'h65, 8'h7B},
{8'h85, 8'h81, 8'h88},
{8'h85, 8'h7C, 8'h7D},
{8'h87, 8'h7A, 8'h7D},
{8'h84, 8'h79, 8'h7A},
{8'h85, 8'h7F, 8'h73},
{8'h82, 8'h81, 8'h6B},
{8'h80, 8'h7B, 8'h7D},
{8'h7D, 8'h7C, 8'h80},
{8'h7D, 8'h7E, 8'h84},
{8'h7D, 8'h7E, 8'h86},
{8'h7D, 8'h7E, 8'h84},
{8'h7D, 8'h7B, 8'h81},
{8'h82, 8'h7C, 8'h7F},
{8'h82, 8'h7A, 8'h7B},
{8'h80, 8'h7C, 8'h7D},
{8'h82, 8'h7F, 8'h80},
{8'h80, 8'h7E, 8'h7E},
{8'h7E, 8'h7E, 8'h7E},
{8'h7D, 8'h7E, 8'h7D},
{8'h7C, 8'h80, 8'h7E},
{8'h79, 8'h7F, 8'h7D},
{8'h79, 8'h7F, 8'h7D},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'h7F, 8'h7C, 8'h83},
{8'h7F, 8'h7C, 8'h83},
{8'h7F, 8'h7C, 8'h84},
{8'h7F, 8'h7C, 8'h84},
{8'h81, 8'h7F, 8'h83},
{8'h7F, 8'h7E, 8'h7B},
{8'h7D, 8'h7D, 8'h73},
{8'hC3, 8'hC4, 8'hB4},
{8'hF5, 8'hFE, 8'hD0},
{8'hEB, 8'hF3, 8'hC1},
{8'hEF, 8'hF8, 8'hC3},
{8'hDA, 8'hE1, 8'hAC},
{8'hB5, 8'hB7, 8'h88},
{8'hC6, 8'hC5, 8'hA0},
{8'hA5, 8'hA2, 8'h85},
{8'hF5, 8'hF3, 8'hDD},
{8'hF9, 8'hFD, 8'hE6},
{8'hFF, 8'hF8, 8'hE2},
{8'hD0, 8'hA3, 8'h8F},
{8'h6B, 8'h2E, 8'h1D},
{8'hAA, 8'h7F, 8'h64},
{8'hFA, 8'hE8, 8'hCD},
{8'hFC, 8'hF1, 8'hDF},
{8'hF9, 8'hEE, 8'hE0},
{8'hFE, 8'hF5, 8'hD1},
{8'hFD, 8'hF8, 8'hE1},
{8'hFD, 8'hFB, 8'hF6},
{8'hF8, 8'hF8, 8'hF4},
{8'hFA, 8'hF7, 8'hED},
{8'hFF, 8'hFD, 8'hF5},
{8'hA9, 8'h9D, 8'hA4},
{8'h24, 8'h16, 8'h2F},
{8'h04, 8'h04, 8'h1F},
{8'h00, 8'h01, 8'h11},
{8'h04, 8'h09, 8'h1A},
{8'h02, 8'h04, 8'h22},
{8'h06, 8'h00, 8'h26},
{8'h06, 8'h01, 8'h1B},
{8'h05, 8'h03, 8'h17},
{8'h07, 8'h08, 8'h1C},
{8'hB4, 8'hA3, 8'hB1},
{8'hEB, 8'hD5, 8'hDD},
{8'hF6, 8'hE6, 8'hE9},
{8'hFF, 8'hF8, 8'hFB},
{8'hFF, 8'hFC, 8'hFF},
{8'hFE, 8'hFE, 8'hFF},
{8'hFF, 8'hFE, 8'hFF},
{8'hFF, 8'hFB, 8'hFD},
{8'hFC, 8'hF8, 8'hF6},
{8'hFC, 8'hF8, 8'hF7},
{8'hFC, 8'hF8, 8'hF8},
{8'hFC, 8'hF8, 8'hFA},
{8'hFF, 8'hFD, 8'hFF},
{8'hFF, 8'hFE, 8'hFF},
{8'hFF, 8'hFF, 8'hFF},
{8'hFF, 8'hFD, 8'hFF},
{8'hE3, 8'hD3, 8'hDA},
{8'hDD, 8'hCC, 8'hD2},
{8'hF7, 8'hEF, 8'hF2},
{8'hFD, 8'hFB, 8'hFA},
{8'hFF, 8'hFE, 8'hFB},
{8'hFF, 8'hFD, 8'hF9},
{8'hFF, 8'hFD, 8'hF7},
{8'hFF, 8'hF9, 8'hF4},
{8'hFF, 8'hF1, 8'hED},
{8'hFE, 8'hF2, 8'hF3},
{8'hFF, 8'hFF, 8'hFF},
{8'hB1, 8'hBF, 8'hD5},
{8'h21, 8'h38, 8'h6E},
{8'h19, 8'h34, 8'h76},
{8'h0C, 8'h24, 8'h69},
{8'h07, 8'h19, 8'h5A},
{8'h10, 8'h0E, 8'h45},
{8'h09, 8'h07, 8'h39},
{8'h04, 8'h08, 8'h36},
{8'h04, 8'h0E, 8'h3A},
{8'h0D, 8'h1D, 8'h4F},
{8'h16, 8'h2E, 8'h6D},
{8'h21, 8'h41, 8'h8D},
{8'h27, 8'h4B, 8'hA1},
{8'h18, 8'h54, 8'hB6},
{8'h17, 8'h56, 8'hB8},
{8'h11, 8'h51, 8'hB5},
{8'h16, 8'h56, 8'hB8},
{8'h17, 8'h55, 8'hB4},
{8'h1D, 8'h57, 8'hB0},
{8'h18, 8'h4B, 8'hA0},
{8'h11, 8'h38, 8'h88},
{8'h06, 8'h27, 8'h5B},
{8'h01, 8'h1F, 8'h50},
{8'h00, 8'h14, 8'h44},
{8'h01, 8'h0D, 8'h3A},
{8'h07, 8'h11, 8'h3A},
{8'h09, 8'h12, 8'h35},
{8'h0C, 8'h13, 8'h30},
{8'h0D, 8'h14, 8'h2F},
{8'h0C, 8'h17, 8'h44},
{8'h0B, 8'h1C, 8'h50},
{8'h0B, 8'h26, 8'h60},
{8'h0C, 8'h2E, 8'h6E},
{8'h14, 8'h3B, 8'h82},
{8'h14, 8'h42, 8'h8E},
{8'h17, 8'h4A, 8'h99},
{8'h14, 8'h46, 8'h9C},
{8'h26, 8'h3E, 8'hC6},
{8'h27, 8'h40, 8'hA6},
{8'h38, 8'h57, 8'h85},
{8'h4D, 8'h6B, 8'h73},
{8'h53, 8'h6D, 8'h6B},
{8'h67, 8'h78, 8'h7C},
{8'h76, 8'h7E, 8'h8A},
{8'h79, 8'h7C, 8'h89},
{8'h82, 8'h7B, 8'h71},
{8'h82, 8'h7F, 8'h75},
{8'h7E, 8'h80, 8'h7C},
{8'h75, 8'h7C, 8'h7C},
{8'h77, 8'h80, 8'h81},
{8'h7C, 8'h83, 8'h82},
{8'h7C, 8'h7F, 8'h7B},
{8'h7A, 8'h79, 8'h73},
{8'h81, 8'h79, 8'h77},
{8'h7A, 8'h74, 8'h71},
{8'h7D, 8'h77, 8'h73},
{8'h7F, 8'h7A, 8'h77},
{8'h80, 8'h7A, 8'h77},
{8'h82, 8'h7C, 8'h79},
{8'h7C, 8'h78, 8'h74},
{8'h7F, 8'h7A, 8'h78},
{8'h80, 8'h7D, 8'h80},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'h7F, 8'h7D, 8'h7E},
{8'hFF, 8'hD7, 8'h00},
{8'h7F, 8'h7C, 8'h82},
{8'h7F, 8'h7C, 8'h84},
{8'h7F, 8'h7D, 8'h82},
{8'h7C, 8'h7A, 8'h7A},
{8'h7B, 8'h7A, 8'h75},
{8'h93, 8'h93, 8'h88},
{8'hCF, 8'hD7, 8'hAF},
{8'hE9, 8'hF3, 8'hC5},
{8'hEC, 8'hF3, 8'hC2},
{8'hF4, 8'hF9, 8'hC6},
{8'hFA, 8'hFB, 8'hCD},
{8'hE1, 8'hDE, 8'hBA},
{8'hEA, 8'hE4, 8'hCD},
{8'hFC, 8'hF7, 8'hE6},
{8'hFA, 8'hFD, 8'hDD},
{8'hF8, 8'hE7, 8'hCF},
{8'h87, 8'h46, 8'h3A},
{8'h49, 8'h04, 8'h00},
{8'h86, 8'h5E, 8'h4B},
{8'hFF, 8'hF9, 8'hDF},
{8'hFD, 8'hF4, 8'hDE},
{8'hF0, 8'hD5, 8'hC1},
{8'hFB, 8'hDE, 8'hAF},
{8'hFF, 8'hF1, 8'hD7},
{8'hFB, 8'hF7, 8'hF3},
{8'hF9, 8'hFA, 8'hF7},
{8'hFD, 8'hF9, 8'hE7},
{8'hFF, 8'hF9, 8'hE2},
{8'h99, 8'h83, 8'h78},
{8'h24, 8'h0D, 8'h15},
{8'h16, 8'h04, 8'h0D},
{8'h45, 8'h43, 8'h3E},
{8'h07, 8'h0D, 8'h13},
{8'h03, 8'h03, 8'h27},
{8'h07, 8'h00, 8'h29},
{8'h09, 8'h01, 8'h17},
{8'h04, 8'h03, 8'h16},
{8'h00, 8'h03, 8'h25},
{8'h71, 8'h6E, 8'h89},
{8'hE8, 8'hD7, 8'hE5},
{8'hED, 8'hD0, 8'hD3},
{8'hF1, 8'hD9, 8'hDC},
{8'hF9, 8'hEB, 8'hF5},
{8'hFA, 8'hF4, 8'hFB},
{8'hF9, 8'hEF, 8'hF5},
{8'hF3, 8'hE0, 8'hE1},
{8'hE9, 8'hD5, 8'hD9},
{8'hE9, 8'hD5, 8'hDA},
{8'hE8, 8'hD5, 8'hDB},
{8'hE7, 8'hD6, 8'hDC},
{8'hEB, 8'hDD, 8'hE3},
{8'hEF, 8'hE3, 8'hE9},
{8'hF6, 8'hEA, 8'hF0},
{8'hFA, 8'hF1, 8'hF6},
{8'hEA, 8'hD0, 8'hD9},
{8'hD5, 8'hBC, 8'hC3},
{8'hE4, 8'hD0, 8'hD5},
{8'hEE, 8'hE1, 8'hE3},
{8'hF3, 8'hE8, 8'hE9},
{8'hF2, 8'hE3, 8'hE4},
{8'hEF, 8'hDE, 8'hDF},
{8'hEF, 8'hD9, 8'hDC},
{8'hF9, 8'hD2, 8'hDD},
{8'hF3, 8'hD2, 8'hD4},
{8'hF1, 8'hE0, 8'hDD},
{8'hC6, 8'hC2, 8'hC9},
{8'h06, 8'h08, 8'h24},
{8'h00, 8'h00, 8'h21},
{8'h00, 8'h00, 8'h1F},
{8'h00, 8'h00, 8'h16},
{8'h00, 8'h08, 8'h30},
{8'h0E, 8'h1D, 8'h51},
{8'h16, 8'h28, 8'h6F},
{8'h20, 8'h3B, 8'h92},
{8'h1F, 8'h42, 8'hA1},
{8'h1B, 8'h47, 8'hA6},
{8'h16, 8'h46, 8'hA1},
{8'h12, 8'h41, 8'h97},
{8'h16, 8'h3D, 8'h88},
{8'h1A, 8'h42, 8'h8E},
{8'h22, 8'h50, 8'hA0},
{8'h21, 8'h52, 8'hA6},
{8'h19, 8'h4B, 8'hA1},
{8'h14, 8'h40, 8'h95},
{8'h0E, 8'h38, 8'h8C},
{8'h15, 8'h39, 8'h8C},
{8'h1E, 8'h37, 8'h91},
{8'h1E, 8'h3C, 8'h98},
{8'h1E, 8'h43, 8'hA1},
{8'h1E, 8'h48, 8'hAA},
{8'h1B, 8'h4B, 8'hB1},
{8'h17, 8'h4D, 8'hB6},
{8'h15, 8'h4F, 8'hBB},
{8'h15, 8'h50, 8'hBD},
{8'h1C, 8'h4D, 8'hB6},
{8'h1A, 8'h4F, 8'hB8},
{8'h14, 8'h52, 8'hBB},
{8'h0F, 8'h56, 8'hBE},
{8'h0B, 8'h5A, 8'hBE},
{8'h0A, 8'h5C, 8'hBB},
{8'h0B, 8'h5F, 8'hB8},
{8'h09, 8'h5A, 8'hB1},
{8'h10, 8'h46, 8'h9B},
{8'h09, 8'h49, 8'h99},
{8'h03, 8'h4C, 8'h99},
{8'h05, 8'h4A, 8'h99},
{8'h15, 8'h4D, 8'h9F},
{8'h2A, 8'h4F, 8'h96},
{8'h2F, 8'h41, 8'h71},
{8'h51, 8'h56, 8'h6D},
{8'hA7, 8'h8D, 8'h74},
{8'h9F, 8'h89, 8'h70},
{8'h7E, 8'h73, 8'h64},
{8'h80, 8'h7E, 8'h76},
{8'h7F, 8'h82, 8'h7D},
{8'h79, 8'h7B, 8'h77},
{8'h7A, 8'h79, 8'h72},
{8'h92, 8'h8F, 8'h86},
{8'hB4, 8'hAD, 8'hA6},
{8'hB8, 8'hAD, 8'hA6},
{8'hA8, 8'h9C, 8'h95},
{8'h9B, 8'h8B, 8'h86},
{8'h94, 8'h81, 8'h7D},
{8'h96, 8'h82, 8'h7E},
{8'h9F, 8'h89, 8'h86},
{8'h8D, 8'h78, 8'h76},
{8'h80, 8'h7C, 8'h7F},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'h7F, 8'h7E, 8'h78},
{8'h7F, 8'h7E, 8'h7A},
{8'hFF, 8'hD7, 8'h00},
{8'h7F, 8'h7D, 8'h82},
{8'h7D, 8'h7B, 8'h81},
{8'h80, 8'h7E, 8'h81},
{8'h7F, 8'h7D, 8'h7D},
{8'h7D, 8'h7D, 8'h78},
{8'h92, 8'h9A, 8'h7C},
{8'hE9, 8'hF0, 8'hCA},
{8'hEB, 8'hF2, 8'hC4},
{8'hEE, 8'hF3, 8'hC1},
{8'hEB, 8'hEC, 8'hC0},
{8'hDE, 8'hD9, 8'hB7},
{8'hFE, 8'hF5, 8'hE0},
{8'hFD, 8'hF6, 8'hE7},
{8'hFF, 8'hFF, 8'hD6},
{8'hC4, 8'h9F, 8'h83},
{8'h79, 8'h30, 8'h29},
{8'h45, 8'h03, 8'h01},
{8'h8E, 8'h69, 8'h5F},
{8'hFF, 8'hFB, 8'hE4},
{8'hFF, 8'hF2, 8'hD8},
{8'hEE, 8'hCB, 8'hB1},
{8'hF0, 8'hC0, 8'h91},
{8'hF8, 8'hE1, 8'hC5},
{8'hFA, 8'hEE, 8'hE4},
{8'hF8, 8'hEA, 8'hD6},
{8'hFE, 8'hE9, 8'hBF},
{8'hFF, 8'hEC, 8'hBE},
{8'hF4, 8'hEA, 8'hD3},
{8'hB3, 8'hA9, 8'hAB},
{8'hA1, 8'h86, 8'h86},
{8'hB5, 8'hAC, 8'h99},
{8'h07, 8'h0D, 8'h0D},
{8'h01, 8'h00, 8'h29},
{8'h09, 8'h00, 8'h2C},
{8'h0C, 8'h01, 8'h14},
{8'h04, 8'h03, 8'h15},
{8'h04, 8'h0F, 8'h39},
{8'h30, 8'h39, 8'h59},
{8'hD0, 8'hC4, 8'hD3},
{8'hEC, 8'hCB, 8'hCE},
{8'hEF, 8'hCD, 8'hD0},
{8'hE3, 8'hCE, 8'hDC},
{8'hE2, 8'hD4, 8'hE6},
{8'hE6, 8'hD0, 8'hD9},
{8'hE8, 8'hC5, 8'hC6},
{8'hEB, 8'hC9, 8'hD4},
{8'hEB, 8'hCA, 8'hD6},
{8'hEA, 8'hCB, 8'hD5},
{8'hE8, 8'hCC, 8'hD4},
{8'hE5, 8'hCB, 8'hD1},
{8'hE3, 8'hCC, 8'hD2},
{8'hE4, 8'hD0, 8'hD2},
{8'hE6, 8'hD1, 8'hD4},
{8'hE5, 8'hC3, 8'hCA},
{8'hD8, 8'hB8, 8'hBE},
{8'hE1, 8'hC7, 8'hCD},
{8'hE7, 8'hD0, 8'hD6},
{8'hE8, 8'hD3, 8'hD8},
{8'hE7, 8'hCF, 8'hD7},
{8'hE6, 8'hCC, 8'hD5},
{8'hE6, 8'hC9, 8'hD5},
{8'hEF, 8'hC6, 8'hDD},
{8'hEB, 8'hCC, 8'hCF},
{8'hED, 8'hDB, 8'hCC},
{8'hBD, 8'hB6, 8'hAA},
{8'h84, 8'h7F, 8'h84},
{8'h4B, 8'h48, 8'h53},
{8'h36, 8'h32, 8'h30},
{8'h29, 8'h26, 8'h1C},
{8'h1B, 8'h1C, 8'h26},
{8'h1A, 8'h1F, 8'h25},
{8'h0F, 8'h15, 8'h17},
{8'h03, 8'h0B, 8'h0F},
{8'h00, 8'h03, 8'h0F},
{8'h00, 8'h02, 8'h18},
{8'h00, 8'h00, 8'h22},
{8'h00, 8'h00, 8'h26},
{8'h00, 8'h00, 8'h17},
{8'h00, 8'h00, 8'h1D},
{8'h00, 8'h0E, 8'h3A},
{8'h15, 8'h31, 8'h6B},
{8'h1F, 8'h4B, 8'h92},
{8'h22, 8'h56, 8'hA6},
{8'h22, 8'h5B, 8'hB0},
{8'h1C, 8'h57, 8'hAF},
{8'h1E, 8'h57, 8'hB2},
{8'h1D, 8'h57, 8'hB2},
{8'h1C, 8'h59, 8'hB1},
{8'h18, 8'h59, 8'hB1},
{8'h12, 8'h56, 8'hAF},
{8'h0F, 8'h57, 8'hB2},
{8'h0D, 8'h58, 8'hB6},
{8'h0E, 8'h59, 8'hB8},
{8'h13, 8'h56, 8'hA4},
{8'h13, 8'h57, 8'hA6},
{8'h12, 8'h5A, 8'hAE},
{8'h11, 8'h5B, 8'hB4},
{8'h13, 8'h5A, 8'hB5},
{8'h11, 8'h53, 8'hAE},
{8'h16, 8'h53, 8'hAB},
{8'h08, 8'h3A, 8'h8D},
{8'h10, 8'h3F, 8'h71},
{8'h19, 8'h5A, 8'h9B},
{8'h0B, 8'h54, 8'hB7},
{8'h0B, 8'h52, 8'hD0},
{8'h17, 8'h4E, 8'hC4},
{8'h30, 8'h4C, 8'h91},
{8'h83, 8'h88, 8'h7D},
{8'hE1, 8'hD3, 8'h90},
{8'hE6, 8'hAF, 8'h82},
{8'h91, 8'h5F, 8'h3D},
{8'h4D, 8'h29, 8'h14},
{8'h79, 8'h62, 8'h57},
{8'h81, 8'h74, 8'h6D},
{8'h93, 8'h87, 8'h83},
{8'hD1, 8'hC8, 8'hC1},
{8'hFA, 8'hF0, 8'hE7},
{8'hFF, 8'hF7, 8'hEA},
{8'hFF, 8'hF8, 8'hEB},
{8'hFF, 8'hF6, 8'hEB},
{8'hFF, 8'hF0, 8'hE6},
{8'hF7, 8'hE3, 8'hDB},
{8'hF3, 8'hD4, 8'hCE},
{8'hCA, 8'hA1, 8'h9B},
{8'h97, 8'h6E, 8'h6B},
{8'h7F, 8'h7B, 8'h7E},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'h7F, 8'h7E, 8'h7B},
{8'h7F, 8'h7E, 8'h7B},
{8'h7F, 8'h7E, 8'h7C},
{8'h7F, 8'h7D, 8'h7F},
{8'h80, 8'h7D, 8'h85},
{8'h82, 8'h80, 8'h86},
{8'h78, 8'h76, 8'h79},
{8'h7E, 8'h7D, 8'h78},
{8'hCA, 8'hD7, 8'hB2},
{8'hEE, 8'hF8, 8'hD0},
{8'hEE, 8'hF2, 8'hCB},
{8'hED, 8'hEC, 8'hC6},
{8'hD7, 8'hD2, 8'hB2},
{8'hF8, 8'hF4, 8'hDB},
{8'hF6, 8'hEF, 8'hDC},
{8'hFD, 8'hF9, 8'hE8},
{8'hF2, 8'hEE, 8'hC2},
{8'hCC, 8'hA6, 8'h88},
{8'h7C, 8'h31, 8'h29},
{8'h46, 8'h02, 8'h03},
{8'hA7, 8'h84, 8'h78},
{8'hFF, 8'hFD, 8'hE5},
{8'hFF, 8'hFC, 8'hE1},
{8'hBF, 8'h98, 8'h7F},
{8'h9A, 8'h59, 8'h36},
{8'hEB, 8'hC2, 8'hAA},
{8'hFD, 8'hF5, 8'hE4},
{8'hEB, 8'hCF, 8'hB5},
{8'hD8, 8'hAA, 8'h7F},
{8'hF2, 8'hC4, 8'h94},
{8'hFD, 8'hE0, 8'hBD},
{8'hFF, 8'hF9, 8'hE3},
{8'hFF, 8'hFC, 8'hDE},
{8'hEA, 8'hE6, 8'hC9},
{8'h4F, 8'h50, 8'h4E},
{8'h01, 8'h00, 8'h21},
{8'h06, 8'h01, 8'h27},
{8'h09, 8'h04, 8'h15},
{8'h03, 8'h02, 8'h18},
{8'h10, 8'h1A, 8'h4B},
{8'h24, 8'h3E, 8'h70},
{8'h8C, 8'h8F, 8'hA9},
{8'hE9, 8'hD0, 8'hD3},
{8'hEE, 8'hC9, 8'hC9},
{8'hE6, 8'hC6, 8'hD2},
{8'hE0, 8'hC9, 8'hDE},
{8'hE1, 8'hCC, 8'hDA},
{8'hE8, 8'hCE, 8'hD3},
{8'hED, 8'hCA, 8'hD7},
{8'hEC, 8'hC9, 8'hD8},
{8'hEB, 8'hCA, 8'hD7},
{8'hE9, 8'hCB, 8'hD5},
{8'hE8, 8'hCB, 8'hD3},
{8'hE7, 8'hCB, 8'hD0},
{8'hE7, 8'hCC, 8'hCF},
{8'hE7, 8'hCC, 8'hCD},
{8'hEE, 8'hCB, 8'hD3},
{8'hE9, 8'hC8, 8'hCF},
{8'hEB, 8'hCD, 8'hD4},
{8'hE5, 8'hCB, 8'hD2},
{8'hE5, 8'hCB, 8'hD3},
{8'hE8, 8'hCD, 8'hD7},
{8'hEA, 8'hCE, 8'hD9},
{8'hE9, 8'hCB, 8'hD9},
{8'hEC, 8'hC9, 8'hE2},
{8'hE6, 8'hC9, 8'hD2},
{8'hE1, 8'hD0, 8'hC6},
{8'hC3, 8'hB9, 8'hAC},
{8'hF4, 8'hED, 8'hE6},
{8'hE6, 8'hE1, 8'hD7},
{8'hD8, 8'hD5, 8'hB9},
{8'hC0, 8'hC0, 8'h92},
{8'hA7, 8'hB8, 8'h89},
{8'hAC, 8'hBC, 8'h95},
{8'hB2, 8'hBD, 8'hA4},
{8'h99, 8'hA0, 8'h96},
{8'hB3, 8'hB5, 8'hB2},
{8'hB5, 8'hB3, 8'hAD},
{8'hA0, 8'h9E, 8'h91},
{8'h84, 8'h80, 8'h71},
{8'h76, 8'h6B, 8'h61},
{8'h54, 8'h4F, 8'h4F},
{8'h39, 8'h39, 8'h47},
{8'h23, 8'h26, 8'h45},
{8'h05, 8'h13, 8'h3F},
{8'h00, 8'h1B, 8'h55},
{8'h0A, 8'h34, 8'h7B},
{8'h19, 8'h45, 8'h96},
{8'h18, 8'h50, 8'hBA},
{8'h18, 8'h52, 8'hBD},
{8'h18, 8'h52, 8'hBB},
{8'h16, 8'h53, 8'hB8},
{8'h15, 8'h54, 8'hB4},
{8'h14, 8'h55, 8'hAF},
{8'h17, 8'h59, 8'hAC},
{8'h15, 8'h58, 8'hAB},
{8'h13, 8'h56, 8'hC1},
{8'h12, 8'h54, 8'hC4},
{8'h10, 8'h54, 8'hC2},
{8'h12, 8'h53, 8'hBF},
{8'h18, 8'h50, 8'hB5},
{8'h26, 8'h53, 8'hAE},
{8'h1D, 8'h3A, 8'h8C},
{8'h0B, 8'h1E, 8'h69},
{8'h26, 8'h4B, 8'h9B},
{8'h1D, 8'h4C, 8'hB9},
{8'h17, 8'h52, 8'hC7},
{8'h1B, 8'h56, 8'hBE},
{8'h2C, 8'h51, 8'h9B},
{8'h94, 8'h9C, 8'h80},
{8'hFA, 8'hE2, 8'h88},
{8'hCB, 8'h96, 8'h37},
{8'h97, 8'h5A, 8'h30},
{8'hC7, 8'h97, 8'h77},
{8'hDA, 8'hC2, 8'hAC},
{8'hD7, 8'hBD, 8'hB1},
{8'hD8, 8'hC4, 8'hBE},
{8'hF8, 8'hE7, 8'hE4},
{8'hFF, 8'hF2, 8'hEF},
{8'hFF, 8'hF0, 8'hEA},
{8'hFF, 8'hF2, 8'hE4},
{8'hFF, 8'hF7, 8'hEA},
{8'hE0, 8'hCF, 8'hC3},
{8'hC5, 8'hB0, 8'hA7},
{8'hBC, 8'hA7, 8'hA0},
{8'hA8, 8'h8C, 8'h88},
{8'h95, 8'h73, 8'h71},
{8'h90, 8'h6F, 8'h6F},
{8'h82, 8'h7C, 8'h7F},
{8'h81, 8'h7C, 8'h80},
{8'h80, 8'h7C, 8'h80},
{8'h7F, 8'h7C, 8'h80},
{8'h80, 8'h7D, 8'h81},
{8'h7F, 8'h7C, 8'h81},
{8'h7F, 8'h7D, 8'h81},
{8'h80, 8'h7E, 8'h82},
{8'h7F, 8'h7C, 8'h88},
{8'hFF, 8'hD7, 8'h00},
{8'h7F, 8'h7E, 8'h79},
{8'h7E, 8'h7D, 8'h7C},
{8'h7D, 8'h7A, 8'h82},
{8'h7E, 8'h7B, 8'h85},
{8'h7D, 8'h7C, 8'h7B},
{8'h82, 8'h84, 8'h73},
{8'hE0, 8'hF1, 8'hB5},
{8'hF1, 8'hFB, 8'hC9},
{8'hF0, 8'hEC, 8'hCD},
{8'hD2, 8'hC2, 8'hB3},
{8'hF5, 8'hE5, 8'hDE},
{8'hFB, 8'hEF, 8'hE5},
{8'hFA, 8'hF8, 8'hE6},
{8'hF4, 8'hF7, 8'hDB},
{8'hD8, 8'hDF, 8'hB1},
{8'hF2, 8'hDC, 8'hB8},
{8'h75, 8'h31, 8'h1D},
{8'h53, 8'h0F, 8'h02},
{8'hBB, 8'h9A, 8'h80},
{8'hFF, 8'hFD, 8'hE0},
{8'hFF, 8'hFC, 8'hE4},
{8'hB0, 8'h87, 8'h78},
{8'h79, 8'h20, 8'h0D},
{8'hD9, 8'hA0, 8'h8C},
{8'hFF, 8'hF5, 8'hE2},
{8'hF4, 8'hE3, 8'hD6},
{8'h9B, 8'h71, 8'h65},
{8'hD0, 8'h9C, 8'h84},
{8'hE9, 8'hB9, 8'h89},
{8'hDF, 8'hC1, 8'h7C},
{8'hEF, 8'hE3, 8'h93},
{8'hFF, 8'hF8, 8'hCE},
{8'hDC, 8'hD6, 8'hD4},
{8'h0D, 8'h0E, 8'h1E},
{8'h00, 8'h05, 8'h14},
{8'h00, 8'h05, 8'h18},
{8'h00, 8'h00, 8'h21},
{8'h14, 8'h16, 8'h4C},
{8'h1A, 8'h4E, 8'hA8},
{8'h36, 8'h5C, 8'h94},
{8'hC7, 8'hCC, 8'hD9},
{8'hE9, 8'hCD, 8'hC9},
{8'hF5, 8'hC7, 8'hCE},
{8'hEF, 8'hC7, 8'hDB},
{8'hDF, 8'hCB, 8'hDE},
{8'hD5, 8'hD0, 8'hD9},
{8'hE6, 8'hCB, 8'hD4},
{8'hE6, 8'hCA, 8'hD5},
{8'hE5, 8'hCB, 8'hD6},
{8'hE5, 8'hCB, 8'hD6},
{8'hE7, 8'hCD, 8'hD7},
{8'hE9, 8'hCC, 8'hD5},
{8'hEA, 8'hCB, 8'hD1},
{8'hEA, 8'hCA, 8'hD0},
{8'hE7, 8'hC8, 8'hD3},
{8'hE7, 8'hC9, 8'hD3},
{8'hE7, 8'hCA, 8'hD4},
{8'hE7, 8'hCC, 8'hD5},
{8'hE7, 8'hCC, 8'hD5},
{8'hE7, 8'hCD, 8'hD6},
{8'hE7, 8'hCD, 8'hD6},
{8'hE5, 8'hCC, 8'hD5},
{8'hE8, 8'hCA, 8'hD4},
{8'hE9, 8'hCC, 8'hD8},
{8'hE2, 8'hCA, 8'hD4},
{8'hC7, 8'hB6, 8'hB8},
{8'hED, 8'hE5, 8'hD8},
{8'hAD, 8'hAD, 8'h90},
{8'hC2, 8'hC9, 8'h9D},
{8'hC5, 8'hD0, 8'h9B},
{8'hDB, 8'hE7, 8'hAF},
{8'hB9, 8'hC2, 8'h95},
{8'hE5, 8'hEA, 8'hD0},
{8'hF2, 8'hF3, 8'hE9},
{8'hFE, 8'hFA, 8'hF8},
{8'hFF, 8'hFC, 8'hFA},
{8'hFE, 8'hF9, 8'hF0},
{8'hFF, 8'hFD, 8'hEF},
{8'hFA, 8'hFF, 8'hEA},
{8'hFA, 8'hFD, 8'hF3},
{8'hF2, 8'hF3, 8'hF4},
{8'hE9, 8'hE8, 8'hEB},
{8'hC5, 8'hC3, 8'hC3},
{8'h65, 8'h63, 8'h66},
{8'h1F, 8'h1A, 8'h2C},
{8'h03, 8'h00, 8'h20},
{8'h03, 8'h10, 8'h47},
{8'h11, 8'h21, 8'h63},
{8'h1D, 8'h39, 8'h89},
{8'h21, 8'h46, 8'hA2},
{8'h20, 8'h51, 8'hB3},
{8'h19, 8'h56, 8'hB4},
{8'h11, 8'h57, 8'hAF},
{8'h0D, 8'h58, 8'hAC},
{8'h0C, 8'h55, 8'hB4},
{8'h0A, 8'h56, 8'hB9},
{8'h09, 8'h57, 8'hBC},
{8'h0B, 8'h57, 8'hBB},
{8'h14, 8'h56, 8'hB3},
{8'h1F, 8'h53, 8'hA6},
{8'h0B, 8'h21, 8'h69},
{8'h11, 8'h20, 8'h60},
{8'h1B, 8'h58, 8'h9D},
{8'h10, 8'h53, 8'hC3},
{8'h10, 8'h54, 8'hC5},
{8'h1F, 8'h51, 8'h98},
{8'h7C, 8'h86, 8'h93},
{8'hFB, 8'hE7, 8'h70},
{8'hCE, 8'h8E, 8'h49},
{8'hA0, 8'h44, 8'h3B},
{8'hDD, 8'hC4, 8'hB1},
{8'hFF, 8'hF9, 8'hE9},
{8'hFF, 8'hF4, 8'hE8},
{8'hFF, 8'hF8, 8'hEF},
{8'hFF, 8'hF6, 8'hF0},
{8'hFD, 8'hF3, 8'hED},
{8'hFD, 8'hF0, 8'hEA},
{8'hFF, 8'hEF, 8'hE8},
{8'hFF, 8'hEB, 8'hE0},
{8'hE7, 8'hD5, 8'hCB},
{8'h9D, 8'h8F, 8'h86},
{8'h74, 8'h6E, 8'h67},
{8'h71, 8'h6F, 8'h6B},
{8'h77, 8'h78, 8'h79},
{8'h7F, 8'h7F, 8'h85},
{8'h7F, 8'h7D, 8'h84},
{8'h84, 8'h7D, 8'h80},
{8'h83, 8'h7D, 8'h7E},
{8'h80, 8'h7A, 8'h7E},
{8'h7E, 8'h79, 8'h7D},
{8'h80, 8'h7C, 8'h82},
{8'h80, 8'h7E, 8'h84},
{8'h7E, 8'h7E, 8'h84},
{8'h7D, 8'h7C, 8'h83},
{8'h7F, 8'h7C, 8'h87},
{8'hFF, 8'hD7, 8'h00},
{8'h7F, 8'h7E, 8'h7A},
{8'h7F, 8'h7D, 8'h7E},
{8'h7D, 8'h7A, 8'h83},
{8'h80, 8'h7C, 8'h86},
{8'h7E, 8'h7D, 8'h79},
{8'h82, 8'h84, 8'h70},
{8'hE2, 8'hE6, 8'hAE},
{8'hF7, 8'hF3, 8'hC4},
{8'hDB, 8'hCC, 8'hAD},
{8'hE5, 8'hD0, 8'hBF},
{8'hFD, 8'hE5, 8'hDA},
{8'hFF, 8'hEE, 8'hE1},
{8'hF6, 8'hEA, 8'hD5},
{8'hDC, 8'hD5, 8'hB8},
{8'hE7, 8'hF3, 8'hBD},
{8'hFC, 8'hEE, 8'hC3},
{8'h8E, 8'h5A, 8'h42},
{8'h5E, 8'h28, 8'h12},
{8'hCF, 8'hB9, 8'h9F},
{8'hFF, 8'hFF, 8'hE5},
{8'hFE, 8'hF4, 8'hDF},
{8'hBF, 8'h9C, 8'h8D},
{8'hAB, 8'h75, 8'h5F},
{8'hCE, 8'hAC, 8'h94},
{8'hF8, 8'hF1, 8'hDB},
{8'hFB, 8'hF3, 8'hE2},
{8'hEB, 8'hD8, 8'hC5},
{8'hFB, 8'hE2, 8'hC5},
{8'hF3, 8'hDC, 8'hAC},
{8'hDE, 8'hD1, 8'h92},
{8'hD2, 8'hBF, 8'h78},
{8'hE3, 8'hD4, 8'hAA},
{8'hB8, 8'hB1, 8'hAB},
{8'h0E, 8'h10, 8'h1D},
{8'h00, 8'h05, 8'h15},
{8'h00, 8'h04, 8'h17},
{8'h00, 8'h01, 8'h21},
{8'h0D, 8'h11, 8'h43},
{8'h12, 8'h50, 8'hB2},
{8'h1C, 8'h50, 8'h99},
{8'h65, 8'h7D, 8'hA1},
{8'hD7, 8'hCE, 8'hE1},
{8'hEE, 8'hCC, 8'hDE},
{8'hF0, 8'hC4, 8'hD5},
{8'hF6, 8'hCB, 8'hCF},
{8'hF2, 8'hCC, 8'hC3},
{8'hE9, 8'hCB, 8'hCE},
{8'hE8, 8'hCB, 8'hD0},
{8'hE7, 8'hCB, 8'hD2},
{8'hE7, 8'hCB, 8'hD2},
{8'hEB, 8'hCF, 8'hD8},
{8'hEC, 8'hCF, 8'hD7},
{8'hEC, 8'hCE, 8'hD6},
{8'hEA, 8'hCC, 8'hD4},
{8'hDC, 8'hC6, 8'hCD},
{8'hE1, 8'hCA, 8'hD2},
{8'hE5, 8'hCE, 8'hD6},
{8'hE5, 8'hCC, 8'hD5},
{8'hE4, 8'hCB, 8'hD4},
{8'hE8, 8'hCE, 8'hD7},
{8'hE9, 8'hCE, 8'hD7},
{8'hE5, 8'hCB, 8'hD3},
{8'hE6, 8'hCC, 8'hCB},
{8'hE7, 8'hCF, 8'hCE},
{8'hD8, 8'hC4, 8'hC1},
{8'hD1, 8'hC3, 8'hBC},
{8'hF0, 8'hE9, 8'hD8},
{8'h9A, 8'h9A, 8'h7D},
{8'hAD, 8'hB2, 8'h8B},
{8'hC7, 8'hCF, 8'hA0},
{8'hC8, 8'hD1, 8'hA7},
{8'hB6, 8'hBD, 8'h9C},
{8'hF6, 8'hF9, 8'hE7},
{8'hF8, 8'hF8, 8'hF1},
{8'hF9, 8'hF6, 8'hF3},
{8'hFA, 8'hF6, 8'hEC},
{8'hE7, 8'hE5, 8'hD1},
{8'hF5, 8'hF4, 8'hDA},
{8'hF4, 8'hF1, 8'hE7},
{8'hF7, 8'hF5, 8'hF3},
{8'hFD, 8'hFB, 8'hFE},
{8'hFF, 8'hFF, 8'hFA},
{8'hFF, 8'hFF, 8'hF3},
{8'hF7, 8'hFC, 8'hE3},
{8'hD4, 8'hDA, 8'hC6},
{8'hA1, 8'hA6, 8'h9C},
{8'h51, 8'h5C, 8'h51},
{8'h14, 8'h1D, 8'h1A},
{8'h00, 8'h06, 8'h16},
{8'h00, 8'h0A, 8'h2F},
{8'h09, 8'h1F, 8'h59},
{8'h11, 8'h2E, 8'h7A},
{8'h19, 8'h3D, 8'h96},
{8'h1F, 8'h45, 8'hA5},
{8'h23, 8'h49, 8'hA4},
{8'h21, 8'h4A, 8'hA6},
{8'h20, 8'h4C, 8'hA7},
{8'h20, 8'h4D, 8'hA4},
{8'h23, 8'h4A, 8'h97},
{8'h1D, 8'h3A, 8'h7B},
{8'h03, 8'h0B, 8'h3F},
{8'h15, 8'h1C, 8'h4D},
{8'h18, 8'h56, 8'hB5},
{8'h0C, 8'h5C, 8'hB6},
{8'h0B, 8'h53, 8'hB7},
{8'h2D, 8'h4E, 8'h94},
{8'hD8, 8'hCF, 8'h8C},
{8'hEC, 8'hBF, 8'h4A},
{8'h92, 8'h45, 8'h2E},
{8'hCA, 8'h94, 8'h78},
{8'hFF, 8'hF8, 8'hE8},
{8'hFC, 8'hF2, 8'hE9},
{8'hFC, 8'hF2, 8'hEA},
{8'hF8, 8'hEF, 8'hE6},
{8'hFA, 8'hEE, 8'hE5},
{8'hF7, 8'hE6, 8'hD9},
{8'hFB, 8'hE7, 8'hD6},
{8'hFF, 8'hF1, 8'hDE},
{8'hFF, 8'hE9, 8'hDD},
{8'hF1, 8'hD9, 8'hCE},
{8'hF4, 8'hE5, 8'hDA},
{8'hE3, 8'hDA, 8'hD1},
{8'hAD, 8'hA4, 8'h9F},
{8'h86, 8'h7C, 8'h7A},
{8'h81, 8'h75, 8'h78},
{8'h82, 8'h78, 8'h7B},
{8'h7F, 8'h7A, 8'h77},
{8'h7E, 8'h7C, 8'h78},
{8'h7F, 8'h7D, 8'h7A},
{8'h7E, 8'h7E, 8'h7C},
{8'h7E, 8'h7F, 8'h7E},
{8'h81, 8'h82, 8'h82},
{8'h7F, 8'h81, 8'h83},
{8'h7B, 8'h7D, 8'h7E},
{8'h7F, 8'h7C, 8'h85},
{8'hFF, 8'hD7, 8'h00},
{8'h7F, 8'h7E, 8'h7B},
{8'hFF, 8'hD7, 8'h00},
{8'h79, 8'h76, 8'h80},
{8'h7E, 8'h7B, 8'h83},
{8'h81, 8'h80, 8'h79},
{8'hB4, 8'hB6, 8'h9D},
{8'hF4, 8'hF0, 8'hBB},
{8'hF7, 8'hED, 8'hBE},
{8'hC3, 8'hAF, 8'h8C},
{8'hF2, 8'hDD, 8'hC4},
{8'hFA, 8'hE2, 8'hCD},
{8'hEA, 8'hD2, 8'hBB},
{8'hE0, 8'hD0, 8'hB3},
{8'hEF, 8'hE6, 8'hC2},
{8'hE5, 8'hFA, 8'hBD},
{8'hFA, 8'hF7, 8'hC3},
{8'hC1, 8'hA3, 8'h80},
{8'hA6, 8'h84, 8'h68},
{8'hDD, 8'hCD, 8'hB2},
{8'hFD, 8'hFA, 8'hE2},
{8'hF9, 8'hF3, 8'hE2},
{8'hE9, 8'hD8, 8'hCD},
{8'hFF, 8'hFC, 8'hE6},
{8'hE0, 8'hD6, 8'hBF},
{8'hF3, 8'hF3, 8'hDE},
{8'hFD, 8'hFD, 8'hEC},
{8'hE4, 8'hE1, 8'hCC},
{8'hF6, 8'hF0, 8'hD2},
{8'hE5, 8'hE2, 8'hB7},
{8'hD5, 8'hD7, 8'hA1},
{8'hE3, 8'hD4, 8'h98},
{8'hF6, 8'hE9, 8'hC2},
{8'hC4, 8'hBD, 8'hB1},
{8'h10, 8'h10, 8'h16},
{8'h00, 8'h04, 8'h11},
{8'h00, 8'h04, 8'h17},
{8'h01, 8'h03, 8'h22},
{8'h06, 8'h0B, 8'h38},
{8'h0E, 8'h4E, 8'hB3},
{8'h19, 8'h58, 8'hB1},
{8'h20, 8'h4D, 8'h90},
{8'h60, 8'h75, 8'hAA},
{8'hBC, 8'hB8, 8'hE1},
{8'hEB, 8'hCE, 8'hE9},
{8'hFA, 8'hCD, 8'hD2},
{8'hFE, 8'hCA, 8'hC1},
{8'hEB, 8'hD0, 8'hD3},
{8'hE9, 8'hD0, 8'hD4},
{8'hE7, 8'hCD, 8'hD2},
{8'hE6, 8'hCB, 8'hD0},
{8'hE7, 8'hCB, 8'hD2},
{8'hE7, 8'hCB, 8'hD4},
{8'hE5, 8'hCA, 8'hD5},
{8'hE2, 8'hC8, 8'hD3},
{8'hD5, 8'hC9, 8'hCD},
{8'hE1, 8'hD5, 8'hD9},
{8'hE9, 8'hDA, 8'hDF},
{8'hE7, 8'hD5, 8'hDC},
{8'hE2, 8'hCC, 8'hD3},
{8'hE7, 8'hCE, 8'hD6},
{8'hEA, 8'hCF, 8'hD8},
{8'hE7, 8'hCB, 8'hD4},
{8'hE7, 8'hD3, 8'hCD},
{8'hE1, 8'hCF, 8'hC8},
{8'hC9, 8'hBA, 8'hB2},
{8'hE6, 8'hDB, 8'hD1},
{8'hF3, 8'hEC, 8'hDC},
{8'hDC, 8'hD9, 8'hC3},
{8'hB1, 8'hB2, 8'h95},
{8'hC6, 8'hC9, 8'hA9},
{8'hC4, 8'hC8, 8'hB0},
{8'hEE, 8'hF0, 8'hDF},
{8'hF7, 8'hF8, 8'hF0},
{8'hF3, 8'hF2, 8'hED},
{8'hF9, 8'hF7, 8'hF0},
{8'hFB, 8'hFA, 8'hE6},
{8'hE3, 8'hE4, 8'hC1},
{8'hDF, 8'hE1, 8'hB7},
{8'hEF, 8'hE8, 8'hDE},
{8'hF4, 8'hED, 8'hED},
{8'hF7, 8'hF3, 8'hF4},
{8'hF9, 8'hF9, 8'hED},
{8'hF6, 8'hFA, 8'hDA},
{8'hE2, 8'hED, 8'hBC},
{8'hE6, 8'hF3, 8'hC0},
{8'hF4, 8'hFE, 8'hD5},
{8'hFF, 8'hFF, 8'hE5},
{8'hD1, 8'hD6, 8'hBB},
{8'h94, 8'h99, 8'h82},
{8'h54, 8'h5A, 8'h4B},
{8'h26, 8'h28, 8'h29},
{8'h00, 8'h04, 8'h18},
{8'h00, 8'h00, 8'h26},
{8'h00, 8'h04, 8'h35},
{8'h01, 8'h04, 8'h3D},
{8'h05, 8'h08, 8'h44},
{8'h06, 8'h0C, 8'h48},
{8'h07, 8'h0E, 8'h48},
{8'h05, 8'h0C, 8'h41},
{8'h03, 8'h06, 8'h33},
{8'h04, 8'h03, 8'h25},
{8'h10, 8'h0F, 8'h30},
{8'h16, 8'h48, 8'hAD},
{8'h0B, 8'h59, 8'hC2},
{8'h08, 8'h58, 8'hB1},
{8'h34, 8'h52, 8'h86},
{8'hF0, 8'hDA, 8'h6E},
{8'hD2, 8'h8D, 8'h2B},
{8'h93, 8'h3D, 8'h39},
{8'hE6, 8'hC5, 8'hA6},
{8'hFE, 8'hFA, 8'hEB},
{8'hFB, 8'hEF, 8'hE6},
{8'hFB, 8'hF2, 8'hE8},
{8'hFE, 8'hF6, 8'hEC},
{8'hFC, 8'hF4, 8'hE8},
{8'hFB, 8'hEC, 8'hDB},
{8'hEF, 8'hD8, 8'hC3},
{8'hDE, 8'hC4, 8'hAE},
{8'hF1, 8'hD4, 8'hC6},
{8'hFF, 8'hE8, 8'hDA},
{8'hFF, 8'hEC, 8'hDF},
{8'hFF, 8'hF5, 8'hE9},
{8'hFF, 8'hF6, 8'hEE},
{8'hF1, 8'hE3, 8'hDE},
{8'hC6, 8'hB4, 8'hB2},
{8'hA6, 8'h91, 8'h90},
{8'h9D, 8'h94, 8'h8D},
{8'h99, 8'h91, 8'h89},
{8'h91, 8'h8B, 8'h83},
{8'h8A, 8'h85, 8'h7E},
{8'h7C, 8'h78, 8'h73},
{8'h7D, 8'h79, 8'h74},
{8'h80, 8'h7E, 8'h7A},
{8'h82, 8'h80, 8'h7D},
{8'h7F, 8'h7C, 8'h84},
{8'h7F, 8'h7D, 8'h7F},
{8'h7F, 8'h7E, 8'h7C},
{8'h7F, 8'h7C, 8'h80},
{8'h80, 8'h7D, 8'h88},
{8'h80, 8'h7D, 8'h83},
{8'h80, 8'h81, 8'h74},
{8'hDE, 8'hE0, 8'hC2},
{8'hF3, 8'hF3, 8'hBF},
{8'hF5, 8'hF1, 8'hC0},
{8'hC7, 8'hBC, 8'h93},
{8'hC3, 8'hB5, 8'h92},
{8'hDA, 8'hCC, 8'hAA},
{8'hE5, 8'hD9, 8'hB5},
{8'hF9, 8'hF4, 8'hCC},
{8'hF0, 8'hF0, 8'hC2},
{8'hE2, 8'hFB, 8'hBB},
{8'hED, 8'hF5, 8'hBC},
{8'hFD, 8'hF3, 8'hC7},
{8'hF7, 8'hE8, 8'hC6},
{8'hED, 8'hE4, 8'hC8},
{8'hFE, 8'hFC, 8'hE6},
{8'hF5, 8'hF0, 8'hE2},
{8'hE1, 8'hD6, 8'hCC},
{8'hFC, 8'hF6, 8'hE4},
{8'hE7, 8'hE0, 8'hCF},
{8'hF7, 8'hF4, 8'hE5},
{8'hFB, 8'hF9, 8'hEB},
{8'hE8, 8'hE6, 8'hD4},
{8'hEE, 8'hED, 8'hD4},
{8'hEF, 8'hF1, 8'hD1},
{8'hE0, 8'hE2, 8'hBC},
{8'hF3, 8'hE6, 8'hB8},
{8'hF4, 8'hE9, 8'hC5},
{8'hF3, 8'hEF, 8'hDA},
{8'h6A, 8'h6A, 8'h65},
{8'h00, 8'h00, 8'h07},
{8'h00, 8'h02, 8'h18},
{8'h05, 8'h06, 8'h23},
{8'h02, 8'h05, 8'h2B},
{8'h0F, 8'h40, 8'h97},
{8'h18, 8'h55, 8'hB0},
{8'h18, 8'h54, 8'hAF},
{8'h1B, 8'h50, 8'hA5},
{8'h29, 8'h4D, 8'h97},
{8'h4F, 8'h5A, 8'h91},
{8'h7E, 8'h71, 8'h93},
{8'h9C, 8'h83, 8'h97},
{8'hAD, 8'hA1, 8'hAF},
{8'hC0, 8'hB3, 8'hBF},
{8'hD6, 8'hC5, 8'hCE},
{8'hE6, 8'hD1, 8'hD8},
{8'hDE, 8'hC7, 8'hCE},
{8'hDD, 8'hC7, 8'hCE},
{8'hDD, 8'hC8, 8'hD2},
{8'hE2, 8'hD0, 8'hDA},
{8'hED, 8'hEA, 8'hEC},
{8'hF9, 8'hF6, 8'hF7},
{8'hFD, 8'hF9, 8'hFB},
{8'hFC, 8'hF5, 8'hF9},
{8'hF1, 8'hE3, 8'hE9},
{8'hE3, 8'hCE, 8'hD5},
{8'hD9, 8'hC0, 8'hC9},
{8'hE9, 8'hD0, 8'hD8},
{8'hEB, 8'hDB, 8'hDE},
{8'hDA, 8'hCC, 8'hCD},
{8'hC8, 8'hBB, 8'hBB},
{8'hF1, 8'hE7, 8'hE3},
{8'hF0, 8'hE8, 8'hDF},
{8'hF6, 8'hF0, 8'hE4},
{8'hE4, 8'hE1, 8'hD1},
{8'hC4, 8'hC1, 8'hB1},
{8'hEB, 8'hEB, 8'hDE},
{8'hFB, 8'hFA, 8'hF3},
{8'hF6, 8'hF5, 8'hF3},
{8'hF7, 8'hF6, 8'hF3},
{8'hFC, 8'hFC, 8'hF1},
{8'hF2, 8'hF4, 8'hD9},
{8'hEB, 8'hF0, 8'hC2},
{8'hE5, 8'hEB, 8'hB4},
{8'hE7, 8'hE0, 8'hCB},
{8'hEF, 8'hE7, 8'hDF},
{8'hEC, 8'hE6, 8'hE3},
{8'hE7, 8'hE6, 8'hDB},
{8'hDF, 8'hE3, 8'hC6},
{8'hE3, 8'hEC, 8'hC2},
{8'hDF, 8'hEC, 8'hBF},
{8'hE6, 8'hEF, 8'hCD},
{8'hF5, 8'hF3, 8'hF0},
{8'hF8, 8'hF7, 8'hED},
{8'hF4, 8'hF7, 8'hDC},
{8'hED, 8'hF4, 8'hCC},
{8'hDD, 8'hE6, 8'hBB},
{8'hBC, 8'hC5, 8'h9E},
{8'h97, 8'h9E, 8'h82},
{8'h5B, 8'h61, 8'h4D},
{8'h3A, 8'h3A, 8'h3A},
{8'h16, 8'h15, 8'h1C},
{8'h00, 8'h00, 8'h0E},
{8'h00, 8'h00, 8'h11},
{8'h00, 8'h00, 8'h19},
{8'h04, 8'h03, 8'h20},
{8'h08, 8'h03, 8'h22},
{8'h05, 8'h02, 8'h1E},
{8'h1E, 8'h33, 8'h84},
{8'h14, 8'h4E, 8'hCB},
{8'h07, 8'h5D, 8'hB7},
{8'h28, 8'h54, 8'h88},
{8'hDB, 8'hC6, 8'h6C},
{8'hD6, 8'h87, 8'h46},
{8'h9D, 8'h43, 8'h40},
{8'hD8, 8'hA5, 8'h8A},
{8'hF8, 8'hDE, 8'hC7},
{8'hFF, 8'hED, 8'hD9},
{8'hFF, 8'hF2, 8'hE2},
{8'hFC, 8'hF0, 8'hE3},
{8'hFC, 8'hF0, 8'hE5},
{8'hFF, 8'hF5, 8'hE9},
{8'hFD, 8'hF2, 8'hE4},
{8'hF4, 8'hE5, 8'hD6},
{8'hE2, 8'hBA, 8'hAA},
{8'hDA, 8'hB2, 8'hA4},
{8'hDB, 8'hBC, 8'hAD},
{8'hE2, 8'hC7, 8'hBA},
{8'hFA, 8'hE2, 8'hD7},
{8'hFF, 8'hF5, 8'hEC},
{8'hFE, 8'hE6, 8'hE0},
{8'hF6, 8'hDA, 8'hD6},
{8'hF8, 8'hE4, 8'hDD},
{8'hF6, 8'hE3, 8'hDB},
{8'hF4, 8'hE4, 8'hDD},
{8'hF2, 8'hE6, 8'hE0},
{8'hE7, 8'hD8, 8'hD2},
{8'hC2, 8'hB2, 8'hAE},
{8'h8F, 8'h7F, 8'h7C},
{8'h85, 8'h75, 8'h72},
{8'h7F, 8'h7D, 8'h82},
{8'h7F, 8'h7D, 8'h7F},
{8'h7F, 8'h7D, 8'h7D},
{8'h7F, 8'h7D, 8'h82},
{8'h80, 8'h7C, 8'h88},
{8'h78, 8'h76, 8'h79},
{8'h9A, 8'h9B, 8'h8A},
{8'hEC, 8'hF0, 8'hCB},
{8'hF0, 8'hF8, 8'hC6},
{8'hEE, 8'hF5, 8'hC4},
{8'hEE, 8'hF3, 8'hC5},
{8'hEB, 8'hEE, 8'hC2},
{8'hED, 8'hF3, 8'hC5},
{8'hEE, 8'hF6, 8'hC5},
{8'hEB, 8'hF5, 8'hC2},
{8'hE7, 8'hF4, 8'hBF},
{8'hE2, 8'hF9, 8'hBB},
{8'hE7, 8'hF5, 8'hBD},
{8'hF4, 8'hF5, 8'hC7},
{8'hDE, 8'hD8, 8'hB4},
{8'hF2, 8'hEC, 8'hD0},
{8'hFF, 8'hFB, 8'hE7},
{8'hF7, 8'hF0, 8'hE2},
{8'hDB, 8'hD3, 8'hC8},
{8'hF0, 8'hEB, 8'hDF},
{8'hE5, 8'hD8, 8'hCD},
{8'hEF, 8'hE1, 8'hD8},
{8'hFF, 8'hF3, 8'hE8},
{8'hF5, 8'hEB, 8'hDB},
{8'hE4, 8'hDE, 8'hCB},
{8'hF3, 8'hED, 8'hD9},
{8'hEF, 8'hE6, 8'hD1},
{8'hE1, 8'hD6, 8'hB6},
{8'hE4, 8'hDC, 8'hB9},
{8'hEB, 8'hE8, 8'hCA},
{8'hD6, 8'hD6, 8'hC7},
{8'h1E, 8'h1F, 8'h26},
{8'h00, 8'h01, 8'h14},
{8'h07, 8'h07, 8'h23},
{8'h01, 8'h01, 8'h20},
{8'h07, 8'h1C, 8'h5A},
{8'h24, 8'h50, 8'hA0},
{8'h17, 8'h52, 8'hB4},
{8'h10, 8'h57, 8'hC0},
{8'h0D, 8'h53, 8'hB4},
{8'h18, 8'h4F, 8'hA2},
{8'h10, 8'h33, 8'h7B},
{8'h00, 8'h0D, 8'h4E},
{8'h06, 8'h0D, 8'h33},
{8'h13, 8'h15, 8'h34},
{8'h1F, 8'h1D, 8'h32},
{8'h78, 8'h6F, 8'h7D},
{8'hDB, 8'hCE, 8'hD7},
{8'hF0, 8'hE3, 8'hE9},
{8'hFA, 8'hEF, 8'hF5},
{8'hFE, 8'hF8, 8'hFD},
{8'hFE, 8'hFF, 8'hFF},
{8'hFD, 8'hFD, 8'hFD},
{8'hFC, 8'hFC, 8'hFD},
{8'hFD, 8'hFB, 8'hFD},
{8'hFF, 8'hFA, 8'hFE},
{8'hFF, 8'hF7, 8'hFC},
{8'hF7, 8'hEB, 8'hF0},
{8'hDD, 8'hCD, 8'hD3},
{8'h96, 8'h8B, 8'h9C},
{8'h9A, 8'h90, 8'h9F},
{8'hE6, 8'hDD, 8'hE4},
{8'hEE, 8'hE5, 8'hE5},
{8'hE9, 8'hE0, 8'hDA},
{8'hF5, 8'hED, 8'hE2},
{8'hFC, 8'hF6, 8'hE9},
{8'hF0, 8'hE9, 8'hDC},
{8'hFE, 8'hFB, 8'hF1},
{8'hF8, 8'hF5, 8'hF0},
{8'hF8, 8'hF4, 8'hF4},
{8'hFB, 8'hF9, 8'hF8},
{8'hF6, 8'hF7, 8'hEC},
{8'hEA, 8'hED, 8'hD1},
{8'hE5, 8'hED, 8'hBC},
{8'hD8, 8'hE1, 8'hA6},
{8'hBA, 8'hB9, 8'h94},
{8'hEC, 8'hE8, 8'hD3},
{8'hF2, 8'hEE, 8'hE7},
{8'hF6, 8'hF4, 8'hEF},
{8'hF0, 8'hF0, 8'hE1},
{8'hE6, 8'hE7, 8'hD0},
{8'hE4, 8'hE8, 8'hD2},
{8'hED, 8'hF1, 8'hE2},
{8'hF9, 8'hFB, 8'hF8},
{8'hF2, 8'hF6, 8'hE9},
{8'hE8, 8'hEE, 8'hD2},
{8'hE3, 8'hEB, 8'hC1},
{8'hEA, 8'hF3, 8'hC1},
{8'hEA, 8'hF5, 8'hC2},
{8'hF9, 8'hFF, 8'hD4},
{8'hEB, 8'hF2, 8'hC9},
{8'hCF, 8'hD6, 8'hA8},
{8'hBB, 8'hC3, 8'h9A},
{8'hA0, 8'hA7, 8'h8C},
{8'h5C, 8'h62, 8'h57},
{8'h1B, 8'h20, 8'h24},
{8'h00, 8'h00, 8'h0F},
{8'h00, 8'h00, 8'h1A},
{8'h04, 8'h03, 8'h21},
{8'h13, 8'h0B, 8'h45},
{8'h18, 8'h3C, 8'h9C},
{8'h0E, 8'h5A, 8'hBD},
{8'h23, 8'h56, 8'hAA},
{8'hB9, 8'hB7, 8'h7A},
{8'hE0, 8'h9F, 8'h6B},
{8'h83, 8'h2C, 8'h3A},
{8'hC0, 8'h82, 8'h67},
{8'hE6, 8'hAE, 8'h8A},
{8'hEF, 8'hC2, 8'hA4},
{8'hFB, 8'hDE, 8'hC6},
{8'hFE, 8'hED, 8'hDC},
{8'hFD, 8'hF2, 8'hE8},
{8'hFA, 8'hF1, 8'hEB},
{8'hFA, 8'hF6, 8'hF1},
{8'hF8, 8'hF4, 8'hEE},
{8'hFE, 8'hE5, 8'hD7},
{8'hEA, 8'hC6, 8'hB7},
{8'hE0, 8'hBE, 8'hAF},
{8'hF7, 8'hDE, 8'hCF},
{8'hFF, 8'hEC, 8'hDF},
{8'hFF, 8'hED, 8'hE2},
{8'hFC, 8'hE7, 8'hDE},
{8'hC5, 8'hA3, 8'h9C},
{8'hA4, 8'h82, 8'h7C},
{8'hAA, 8'h89, 8'h84},
{8'hB3, 8'h95, 8'h90},
{8'hC1, 8'hA5, 8'hA2},
{8'hDC, 8'hC1, 8'hBE},
{8'hE8, 8'hD0, 8'hCD},
{8'hD2, 8'hB7, 8'hB5},
{8'h92, 8'h78, 8'h77},
{8'h7F, 8'h7D, 8'h82},
{8'h7F, 8'h7D, 8'h7E},
{8'h7F, 8'h7D, 8'h7F},
{8'h7F, 8'h7C, 8'h84},
{8'h7C, 8'h78, 8'h85},
{8'h7C, 8'h7A, 8'h7C},
{8'hB0, 8'hB2, 8'h9D},
{8'hF5, 8'hFA, 8'hD0},
{8'hEA, 8'hF3, 8'hC7},
{8'hE9, 8'hF3, 8'hC7},
{8'hE9, 8'hF5, 8'hC6},
{8'hE9, 8'hF7, 8'hC5},
{8'hE4, 8'hF4, 8'hC0},
{8'hE1, 8'hF4, 8'hBD},
{8'hE3, 8'hF6, 8'hBE},
{8'hE7, 8'hF9, 8'hC1},
{8'hE8, 8'hF6, 8'hC2},
{8'hE4, 8'hF1, 8'hC0},
{8'hEC, 8'hF4, 8'hC9},
{8'hDA, 8'hD8, 8'hB5},
{8'hF7, 8'hED, 8'hD3},
{8'hFF, 8'hF2, 8'hE0},
{8'hF4, 8'hE7, 8'hD8},
{8'hD8, 8'hD1, 8'hC2},
{8'hEA, 8'hED, 8'hE2},
{8'hC5, 8'hB5, 8'hAD},
{8'hEB, 8'hD4, 8'hCD},
{8'hFF, 8'hED, 8'hE1},
{8'hF8, 8'hE9, 8'hD8},
{8'hDF, 8'hD8, 8'hC5},
{8'hF6, 8'hEA, 8'hDD},
{8'hF8, 8'hE6, 8'hDD},
{8'hDB, 8'hD2, 8'hBE},
{8'hDD, 8'hD8, 8'hB8},
{8'hE0, 8'hDE, 8'hB8},
{8'hF8, 8'hF7, 8'hE0},
{8'h9A, 8'h98, 8'h9C},
{8'h04, 8'h04, 8'h15},
{8'h02, 8'h02, 8'h1D},
{8'h01, 8'h02, 8'h17},
{8'h00, 8'h03, 8'h25},
{8'h18, 8'h2D, 8'h6D},
{8'h24, 8'h53, 8'hB0},
{8'h10, 8'h56, 8'hC1},
{8'h06, 8'h58, 8'hBC},
{8'h05, 8'h53, 8'hAE},
{8'h18, 8'h5A, 8'hB5},
{8'h19, 8'h4E, 8'hAD},
{8'h17, 8'h3D, 8'h81},
{8'h0F, 8'h29, 8'h62},
{8'h08, 8'h11, 8'h3D},
{8'h19, 8'h1D, 8'h36},
{8'hBE, 8'hBD, 8'hCA},
{8'hD0, 8'hCF, 8'hD2},
{8'hB5, 8'hB3, 8'hB3},
{8'hB3, 8'hB2, 8'hB2},
{8'hAE, 8'hAF, 8'hAE},
{8'hA8, 8'hA9, 8'hA9},
{8'hA7, 8'hA6, 8'hA6},
{8'hA9, 8'hA7, 8'hA8},
{8'hB2, 8'hAF, 8'hB0},
{8'hBC, 8'hB7, 8'hB9},
{8'hBB, 8'hB6, 8'hB8},
{8'h97, 8'h90, 8'h95},
{8'h0A, 8'h03, 8'h1C},
{8'h2C, 8'h27, 8'h39},
{8'hF4, 8'hF0, 8'hF5},
{8'hEA, 8'hE4, 8'hDC},
{8'hE6, 8'hE0, 8'hCC},
{8'hEA, 8'hE5, 8'hC8},
{8'hED, 8'hE6, 8'hC6},
{8'hF7, 8'hF1, 8'hD0},
{8'hF9, 8'hF4, 8'hE5},
{8'hF8, 8'hF4, 8'hEB},
{8'hFD, 8'hFA, 8'hF6},
{8'hFE, 8'hFE, 8'hFB},
{8'hE9, 8'hE9, 8'hDF},
{8'hD9, 8'hDD, 8'hC3},
{8'hE7, 8'hF0, 8'hC4},
{8'hB5, 8'hBF, 8'h89},
{8'hAA, 8'hB1, 8'h84},
{8'hD4, 8'hD6, 8'hBB},
{8'hF6, 8'hF5, 8'hEB},
{8'hF9, 8'hF7, 8'hF2},
{8'hFC, 8'hF8, 8'hEC},
{8'hF5, 8'hF2, 8'hDE},
{8'hF0, 8'hEB, 8'hD9},
{8'hED, 8'hE8, 8'hD9},
{8'hE1, 8'hE7, 8'hC6},
{8'hE3, 8'hE9, 8'hC6},
{8'hE5, 8'hEC, 8'hCA},
{8'hE8, 8'hEE, 8'hCD},
{8'hE9, 8'hF0, 8'hD0},
{8'hEF, 8'hF6, 8'hD9},
{8'hF4, 8'hFB, 8'hE1},
{8'hDC, 8'hE4, 8'hCA},
{8'hC4, 8'hD2, 8'h98},
{8'hCF, 8'hDC, 8'hA6},
{8'hDA, 8'hE7, 8'hBB},
{8'hD5, 8'hE0, 8'hC1},
{8'hB2, 8'hBD, 8'hAE},
{8'h89, 8'h91, 8'h91},
{8'h35, 8'h39, 8'h44},
{8'h01, 8'h03, 8'h14},
{8'h0B, 8'h00, 8'h1B},
{8'h03, 8'h14, 8'h3F},
{8'h0F, 8'h40, 8'h99},
{8'h20, 8'h46, 8'hA6},
{8'h95, 8'h9D, 8'h73},
{8'hE6, 8'hC4, 8'h7E},
{8'h3C, 8'h09, 8'h11},
{8'h3F, 8'h12, 8'h0D},
{8'h78, 8'h3B, 8'h23},
{8'hA3, 8'h69, 8'h50},
{8'hCB, 8'h9C, 8'h87},
{8'hE1, 8'hC1, 8'hB2},
{8'hF7, 8'hE2, 8'hD7},
{8'hFF, 8'hF2, 8'hEB},
{8'hFD, 8'hF4, 8'hEC},
{8'hFB, 8'hF1, 8'hE9},
{8'hFF, 8'hE9, 8'hDD},
{8'hFF, 8'hEE, 8'hDF},
{8'hFF, 8'hEF, 8'hE0},
{8'hFE, 8'hEE, 8'hDF},
{8'hF2, 8'hE2, 8'hD4},
{8'hED, 8'hD6, 8'hC9},
{8'hEC, 8'hD8, 8'hCE},
{8'hE0, 8'hC9, 8'hBF},
{8'hBC, 8'hA2, 8'h9B},
{8'h99, 8'h7D, 8'h77},
{8'h85, 8'h6A, 8'h64},
{8'h8A, 8'h70, 8'h6B},
{8'h8B, 8'h72, 8'h6E},
{8'h8D, 8'h75, 8'h71},
{8'h86, 8'h6F, 8'h6D},
{8'h87, 8'h70, 8'h6E},
{8'h7F, 8'h7D, 8'h81},
{8'h7F, 8'h7D, 8'h7E},
{8'h7F, 8'h7D, 8'h7F},
{8'h80, 8'h7C, 8'h86},
{8'h80, 8'h7C, 8'h8A},
{8'h79, 8'h77, 8'h79},
{8'hA8, 8'hAA, 8'h90},
{8'hF1, 8'hF7, 8'hC8},
{8'hEA, 8'hEB, 8'hC8},
{8'hED, 8'hF0, 8'hCB},
{8'hED, 8'hF5, 8'hCA},
{8'hEB, 8'hF8, 8'hC6},
{8'hEA, 8'hF9, 8'hC3},
{8'hED, 8'hFE, 8'hC7},
{8'hEA, 8'hFB, 8'hC4},
{8'hE5, 8'hF4, 8'hBE},
{8'hEF, 8'hF4, 8'hC9},
{8'hE5, 8'hEF, 8'hC4},
{8'hDF, 8'hEA, 8'hC1},
{8'hD3, 8'hD3, 8'hB2},
{8'hFB, 8'hED, 8'hD3},
{8'hFF, 8'hEE, 8'hDC},
{8'hEA, 8'hD8, 8'hC6},
{8'hE5, 8'hDB, 8'hC8},
{8'hDC, 8'hE8, 8'hDC},
{8'hBB, 8'hAF, 8'hA6},
{8'hF3, 8'hDA, 8'hD1},
{8'hFF, 8'hE9, 8'hDB},
{8'hF1, 8'hE0, 8'hCB},
{8'hE0, 8'hDD, 8'hC8},
{8'hF8, 8'hF0, 8'hE3},
{8'hF3, 8'hE1, 8'hDC},
{8'hEC, 8'hE4, 8'hD9},
{8'hD8, 8'hD5, 8'hB6},
{8'hC1, 8'hC0, 8'h94},
{8'hDE, 8'hDD, 8'hBF},
{8'hEF, 8'hED, 8'hEE},
{8'h3E, 8'h3D, 8'h57},
{8'h00, 8'h00, 8'h18},
{8'h01, 8'h03, 8'h13},
{8'h06, 8'h02, 8'h12},
{8'h02, 8'h07, 8'h38},
{8'h1E, 8'h3E, 8'h94},
{8'h14, 8'h4F, 8'hB0},
{8'h0D, 8'h58, 8'hAE},
{8'h0F, 8'h5C, 8'hAA},
{8'h0F, 8'h54, 8'hAC},
{8'h14, 8'h51, 8'hB6},
{8'h1A, 8'h57, 8'hB4},
{8'h21, 8'h55, 8'hA6},
{8'h39, 8'h5E, 8'h9C},
{8'h1D, 8'h31, 8'h56},
{8'h5F, 8'h66, 8'h76},
{8'hBD, 8'hC0, 8'hC2},
{8'hCA, 8'hCE, 8'hCC},
{8'hDE, 8'hE1, 8'hDC},
{8'hEE, 8'hED, 8'hED},
{8'hF5, 8'hF4, 8'hF5},
{8'hF8, 8'hF7, 8'hF8},
{8'hF5, 8'hF5, 8'hF5},
{8'hEF, 8'hEF, 8'hEF},
{8'hE2, 8'hE3, 8'hE2},
{8'hD1, 8'hD2, 8'hD2},
{8'hB1, 8'hB2, 8'hB4},
{8'h2A, 8'h28, 8'h3E},
{8'h3C, 8'h39, 8'h47},
{8'hC7, 8'hC6, 8'hC1},
{8'hE5, 8'hE4, 8'hCA},
{8'hE7, 8'hE5, 8'hB9},
{8'hE1, 8'hDF, 8'hA7},
{8'hD5, 8'hD1, 8'h93},
{8'hEA, 8'hE6, 8'hA7},
{8'hEA, 8'hE5, 8'hCC},
{8'hF3, 8'hEE, 8'hDE},
{8'hFD, 8'hFC, 8'hF3},
{8'hDE, 8'hDB, 8'hD8},
{8'h9D, 8'h9D, 8'h95},
{8'h8D, 8'h91, 8'h7C},
{8'hD1, 8'hD9, 8'hB4},
{8'hB4, 8'hBF, 8'h8F},
{8'hAA, 8'hB6, 8'h89},
{8'hBA, 8'hC3, 8'hA7},
{8'hDF, 8'hE1, 8'hD6},
{8'hF4, 8'hF2, 8'hE9},
{8'hFE, 8'hFB, 8'hE6},
{8'hFE, 8'hFB, 8'hDC},
{8'hFC, 8'hF5, 8'hD1},
{8'hF2, 8'hEA, 8'hC4},
{8'hE6, 8'hE7, 8'hB9},
{8'hEA, 8'hEA, 8'hC4},
{8'hF0, 8'hF0, 8'hD3},
{8'hF4, 8'hF3, 8'hDF},
{8'hF6, 8'hF7, 8'hE7},
{8'hFD, 8'hFE, 8'hEC},
{8'hF2, 8'hF4, 8'hDE},
{8'hE7, 8'hEC, 8'hD1},
{8'hDC, 8'hE8, 8'hC2},
{8'hAD, 8'hB9, 8'h93},
{8'hBE, 8'hC6, 8'hA3},
{8'hBB, 8'hC2, 8'hA2},
{8'hB1, 8'hB7, 8'h9C},
{8'hB3, 8'hBA, 8'hA5},
{8'hC1, 8'hC9, 8'hB8},
{8'h5F, 8'h66, 8'h58},
{8'h02, 8'h05, 8'h01},
{8'h00, 8'h02, 8'h20},
{8'h00, 8'h0A, 8'h47},
{8'h1A, 8'h27, 8'h59},
{8'h7F, 8'h7C, 8'h70},
{8'hE4, 8'hDC, 8'h77},
{8'h3B, 8'h27, 8'h0D},
{8'h12, 8'h00, 8'h08},
{8'h45, 8'h14, 8'h0C},
{8'h66, 8'h36, 8'h2D},
{8'h98, 8'h6D, 8'h63},
{8'hA6, 8'h7E, 8'h73},
{8'hC1, 8'h9C, 8'h8D},
{8'hE5, 8'hC3, 8'hAF},
{8'hFB, 8'hDD, 8'hC6},
{8'hFF, 8'hEB, 8'hD2},
{8'hFB, 8'hE4, 8'hD8},
{8'hF9, 8'hE6, 8'hDA},
{8'hFB, 8'hE9, 8'hDC},
{8'hED, 8'hDA, 8'hCC},
{8'hF1, 8'hE4, 8'hD6},
{8'hFB, 8'hEE, 8'hE0},
{8'hFC, 8'hEB, 8'hDF},
{8'hF5, 8'hE4, 8'hD9},
{8'hE1, 8'hD7, 8'hCC},
{8'hDC, 8'hD0, 8'hC6},
{8'hB6, 8'hAB, 8'hA2},
{8'h89, 8'h80, 8'h77},
{8'h83, 8'h7A, 8'h74},
{8'h82, 8'h7B, 8'h75},
{8'h85, 8'h7E, 8'h78},
{8'h89, 8'h82, 8'h7D},
{8'h7F, 8'h7D, 8'h7F},
{8'h7F, 8'h7D, 8'h7E},
{8'h7F, 8'h7D, 8'h7F},
{8'h7E, 8'h7B, 8'h82},
{8'h81, 8'h7E, 8'h87},
{8'h80, 8'h7E, 8'h7F},
{8'h84, 8'h86, 8'h75},
{8'hD5, 8'hD8, 8'hB9},
{8'hAC, 8'hAB, 8'h8D},
{8'h91, 8'h90, 8'h77},
{8'h98, 8'h9A, 8'h85},
{8'hA2, 8'hA7, 8'h8D},
{8'hAA, 8'hB1, 8'h8E},
{8'hCB, 8'hD5, 8'hA6},
{8'hEE, 8'hF8, 8'hC4},
{8'hEA, 8'hF4, 8'hBD},
{8'hEC, 8'hEF, 8'hC8},
{8'hF0, 8'hF3, 8'hD0},
{8'hE3, 8'hE2, 8'hC4},
{8'hD0, 8'hC3, 8'hA9},
{8'hFD, 8'hE8, 8'hD1},
{8'hFA, 8'hE5, 8'hD3},
{8'hDA, 8'hCB, 8'hBD},
{8'hF1, 8'hE6, 8'hDA},
{8'hCD, 8'hD7, 8'hC2},
{8'hC7, 8'hBD, 8'hAD},
{8'hE8, 8'hCE, 8'hC1},
{8'hFD, 8'hE3, 8'hD2},
{8'hE5, 8'hD3, 8'hBC},
{8'hE9, 8'hE5, 8'hD1},
{8'hF8, 8'hF2, 8'hEA},
{8'hF3, 8'hE7, 8'hE8},
{8'hEB, 8'hE4, 8'hE2},
{8'hD6, 8'hD1, 8'hC0},
{8'hBF, 8'hBC, 8'h9C},
{8'hAD, 8'hAB, 8'h8E},
{8'hDF, 8'hDD, 8'hD2},
{8'hBA, 8'hB7, 8'hBF},
{8'h0A, 8'h08, 8'h1E},
{8'h03, 8'h02, 8'h18},
{8'h0C, 8'h04, 8'h15},
{8'h04, 8'h00, 8'h21},
{8'h09, 8'h13, 8'h52},
{8'h22, 8'h4C, 8'h9B},
{8'h19, 8'h5A, 8'hAC},
{8'h13, 8'h5B, 8'hAF},
{8'h13, 8'h53, 8'hAC},
{8'h19, 8'h4F, 8'hB1},
{8'h12, 8'h53, 8'hBD},
{8'h1F, 8'h55, 8'hAF},
{8'h67, 8'h84, 8'hBF},
{8'h4C, 8'h5E, 8'h86},
{8'h53, 8'h62, 8'h7F},
{8'hF3, 8'hF5, 8'hFA},
{8'hFF, 8'hFF, 8'hFF},
{8'hFC, 8'hFF, 8'hFF},
{8'hFF, 8'hFF, 8'hFF},
{8'hFF, 8'hFF, 8'hFF},
{8'hFE, 8'hFD, 8'hFE},
{8'hFD, 8'hFD, 8'hFD},
{8'hFB, 8'hFC, 8'hFC},
{8'hFB, 8'hFC, 8'hFC},
{8'hFF, 8'hFF, 8'hFF},
{8'hFE, 8'hFF, 8'hFF},
{8'h6E, 8'h6E, 8'h80},
{8'h57, 8'h56, 8'h5F},
{8'h98, 8'h98, 8'h8B},
{8'hF1, 8'hF1, 8'hCD},
{8'hE2, 8'hE1, 8'hA9},
{8'hD4, 8'hD3, 8'h8B},
{8'hBB, 8'hB8, 8'h68},
{8'hDA, 8'hD7, 8'h87},
{8'hEE, 8'hEA, 8'hC9},
{8'hF3, 8'hEE, 8'hDC},
{8'hF7, 8'hF2, 8'hEC},
{8'hF0, 8'hEB, 8'hEB},
{8'hD7, 8'hD5, 8'hD1},
{8'hC8, 8'hC8, 8'hBC},
{8'hD1, 8'hD5, 8'hC1},
{8'hB3, 8'hBA, 8'hA1},
{8'hBF, 8'hC9, 8'hAA},
{8'hBA, 8'hC0, 8'hA6},
{8'hC8, 8'hC8, 8'hB8},
{8'hF9, 8'hF3, 8'hE0},
{8'hF9, 8'hF3, 8'hC1},
{8'hEA, 8'hE3, 8'h90},
{8'hEB, 8'hDE, 8'h8B},
{8'hF8, 8'hEA, 8'hAB},
{8'hF2, 8'hED, 8'hBE},
{8'hF4, 8'hEF, 8'hCA},
{8'hF5, 8'hEF, 8'hD8},
{8'hF4, 8'hEF, 8'hE2},
{8'hFB, 8'hF9, 8'hED},
{8'hF7, 8'hF8, 8'hE2},
{8'hEA, 8'hF1, 8'hCC},
{8'hE5, 8'hEE, 8'hC1},
{8'hEB, 8'hF6, 8'hD2},
{8'hBF, 8'hC8, 8'hA7},
{8'hA7, 8'hAF, 8'h8F},
{8'hC5, 8'hCA, 8'hAF},
{8'hA4, 8'hA8, 8'h90},
{8'h6F, 8'h73, 8'h5E},
{8'h7E, 8'h84, 8'h70},
{8'h92, 8'h99, 8'h85},
{8'h5C, 8'h69, 8'h50},
{8'h0B, 8'h0E, 8'h1B},
{8'h00, 8'h01, 8'h15},
{8'h05, 8'h05, 8'h15},
{8'h43, 8'h38, 8'h43},
{8'hDE, 8'hD9, 8'h7A},
{8'h5D, 8'h51, 8'h1E},
{8'h1C, 8'h04, 8'h1B},
{8'h3C, 8'h19, 8'h1A},
{8'h74, 8'h54, 8'h53},
{8'h95, 8'h79, 8'h79},
{8'h91, 8'h78, 8'h76},
{8'h8F, 8'h74, 8'h6D},
{8'h95, 8'h73, 8'h64},
{8'hB4, 8'h8B, 8'h75},
{8'hCF, 8'hA6, 8'h8D},
{8'hE2, 8'hBF, 8'hAF},
{8'hF9, 8'hDB, 8'hCC},
{8'hFF, 8'hE8, 8'hD8},
{8'hFD, 8'hE7, 8'hD6},
{8'hEA, 8'hCD, 8'hBC},
{8'hD4, 8'hB6, 8'hA6},
{8'hD3, 8'hBA, 8'hA9},
{8'hE2, 8'hCC, 8'hBD},
{8'hD4, 8'hD0, 8'hC4},
{8'hE9, 8'hE4, 8'hD9},
{8'hF6, 8'hF0, 8'hE3},
{8'hE6, 8'hE2, 8'hD5},
{8'hA8, 8'hA5, 8'h99},
{8'h7C, 8'h7A, 8'h72},
{8'h7B, 8'h7F, 8'h7A},
{8'h7C, 8'h81, 8'h7E},
{8'h7F, 8'h7D, 8'h7E},
{8'h7F, 8'h7D, 8'h7E},
{8'h7F, 8'h7D, 8'h7E},
{8'h7F, 8'h7D, 8'h7E},
{8'h7F, 8'h7D, 8'h7D},
{8'h7E, 8'h7C, 8'h7C},
{8'h7B, 8'h79, 8'h7B},
{8'h82, 8'h80, 8'h81},
{8'h85, 8'h89, 8'h70},
{8'h77, 8'h79, 8'h71},
{8'h78, 8'h76, 8'h83},
{8'h76, 8'h74, 8'h81},
{8'h80, 8'h81, 8'h79},
{8'hCC, 8'hD2, 8'hAE},
{8'hEF, 8'hF7, 8'hC2},
{8'hEA, 8'hF4, 8'hB9},
{8'hEB, 8'hF2, 8'hCA},
{8'hF0, 8'hEC, 8'hD3},
{8'hF2, 8'hE6, 8'hDA},
{8'hCD, 8'hAE, 8'hA3},
{8'hFB, 8'hDC, 8'hCC},
{8'hE5, 8'hCD, 8'hBD},
{8'hE6, 8'hDA, 8'hD6},
{8'hFD, 8'hF7, 8'hFB},
{8'hE4, 8'hDE, 8'hBD},
{8'hE3, 8'hD6, 8'hBC},
{8'hD5, 8'hC0, 8'hB1},
{8'hD7, 8'hBE, 8'hAE},
{8'hDF, 8'hC9, 8'hB3},
{8'hFD, 8'hF7, 8'hE4},
{8'hFB, 8'hF6, 8'hF4},
{8'hF3, 8'hF3, 8'hFB},
{8'hE7, 8'hE2, 8'hE3},
{8'hBC, 8'hB6, 8'hB4},
{8'hBC, 8'hB7, 8'hAD},
{8'hA1, 8'hA0, 8'h85},
{8'hD0, 8'hD0, 8'hAC},
{8'hE5, 8'hE2, 8'hCB},
{8'h71, 8'h6A, 8'h72},
{8'h02, 8'h00, 8'h19},
{8'h05, 8'h00, 8'h1B},
{8'h09, 8'h00, 8'h15},
{8'h05, 8'h00, 8'h1D},
{8'h0C, 8'h1C, 8'h53},
{8'h1A, 8'h51, 8'hA9},
{8'h0B, 8'h55, 8'hBF},
{8'h10, 8'h52, 8'hB9},
{8'h1D, 8'h51, 8'hAF},
{8'h19, 8'h51, 8'hBC},
{8'h1F, 8'h4F, 8'hA8},
{8'h54, 8'h63, 8'h96},
{8'h45, 8'h56, 8'h87},
{8'h18, 8'h33, 8'h72},
{8'h8F, 8'h87, 8'h9D},
{8'hCC, 8'hC1, 8'hB3},
{8'hC2, 8'hD5, 8'hD8},
{8'hDA, 8'hE1, 8'hE1},
{8'hE8, 8'hEB, 8'hE9},
{8'hF6, 8'hF6, 8'hF6},
{8'hFF, 8'hFF, 8'hFF},
{8'hFF, 8'hFF, 8'hFF},
{8'hF7, 8'hF2, 8'hF4},
{8'hDB, 8'hD3, 8'hD6},
{8'hC7, 8'hC3, 8'hC6},
{8'h55, 8'h52, 8'h69},
{8'h26, 8'h25, 8'h30},
{8'h6F, 8'h6D, 8'h67},
{8'hEE, 8'hEB, 8'hCE},
{8'hDD, 8'hDA, 8'hAA},
{8'hE5, 8'hE2, 8'hA4},
{8'hCC, 8'hC7, 8'h80},
{8'hDD, 8'hD6, 8'h90},
{8'hE7, 8'hE2, 8'hBF},
{8'hEF, 8'hEA, 8'hD9},
{8'hFA, 8'hF1, 8'hF2},
{8'hF9, 8'hF2, 8'hF7},
{8'hF9, 8'hF4, 8'hF2},
{8'hFC, 8'hF8, 8'hF2},
{8'hF5, 8'hF2, 8'hF2},
{8'hEC, 8'hE9, 8'hEF},
{8'hE3, 8'hE3, 8'hD9},
{8'hC3, 8'hC2, 8'hA8},
{8'hEA, 8'hE4, 8'hCC},
{8'hEF, 8'hE2, 8'hC3},
{8'hE0, 8'hD5, 8'h80},
{8'hDE, 8'hD5, 8'h44},
{8'hEA, 8'hD9, 8'h58},
{8'hF8, 8'hE1, 8'h99},
{8'hF8, 8'hF4, 8'hC0},
{8'hF6, 8'hF3, 8'hC9},
{8'hF7, 8'hF4, 8'hDA},
{8'hFA, 8'hF7, 8'hE9},
{8'hFC, 8'hFC, 8'hEE},
{8'hEE, 8'hF4, 8'hDA},
{8'hE4, 8'hF1, 8'hC4},
{8'hE2, 8'hF2, 8'hB9},
{8'hE7, 8'hF5, 8'hBA},
{8'hE3, 8'hF0, 8'hBC},
{8'hA3, 8'hAE, 8'h87},
{8'hC0, 8'hC9, 8'hAE},
{8'hB9, 8'hC0, 8'hB0},
{8'h7C, 8'h82, 8'h7A},
{8'h81, 8'h86, 8'h81},
{8'h8D, 8'h92, 8'h8F},
{8'hE1, 8'hE4, 8'hD1},
{8'hAA, 8'hB5, 8'h84},
{8'h24, 8'h2F, 8'h18},
{8'h00, 8'h00, 8'h10},
{8'h09, 8'h00, 8'h0B},
{8'h90, 8'h77, 8'h43},
{8'h89, 8'h5B, 8'h30},
{8'h4A, 8'h08, 8'h0B},
{8'h41, 8'h27, 8'h22},
{8'h7C, 8'h6D, 8'h6A},
{8'h82, 8'h7B, 8'h81},
{8'h7E, 8'h7E, 8'h88},
{8'h7B, 8'h7B, 8'h85},
{8'h81, 8'h7A, 8'h80},
{8'h87, 8'h77, 8'h76},
{8'h89, 8'h72, 8'h6B},
{8'hA5, 8'h7A, 8'h6B},
{8'hC3, 8'h98, 8'h88},
{8'hC7, 8'h9D, 8'h8D},
{8'hAE, 8'h85, 8'h75},
{8'h97, 8'h69, 8'h59},
{8'hA4, 8'h76, 8'h66},
{8'hCA, 8'hA0, 8'h90},
{8'hE6, 8'hC2, 8'hB2},
{8'hF4, 8'hE2, 8'hDD},
{8'hF9, 8'hE4, 8'hDC},
{8'hF3, 8'hDA, 8'hCC},
{8'hFA, 8'hDE, 8'hCD},
{8'hFF, 8'hEE, 8'hDF},
{8'hD7, 8'hBD, 8'hB5},
{8'h8C, 8'h7C, 8'h7C},
{8'h82, 8'h78, 8'h7D},
{8'h7F, 8'h7D, 8'h7E},
{8'h7F, 8'h7D, 8'h7E},
{8'h7F, 8'h7D, 8'h7E},
{8'h7F, 8'h7D, 8'h7E},
{8'h7D, 8'h7B, 8'h7C},
{8'h7E, 8'h7C, 8'h7D},
{8'h89, 8'h87, 8'h89},
{8'h83, 8'h82, 8'h81},
{8'h89, 8'h8B, 8'h7F},
{8'h95, 8'h96, 8'h94},
{8'h96, 8'h95, 8'h9A},
{8'hA2, 8'hA2, 8'h9E},
{8'hC3, 8'hC7, 8'hAE},
{8'hF1, 8'hF6, 8'hCA},
{8'hF1, 8'hF8, 8'hC5},
{8'hEA, 8'hF4, 8'hC0},
{8'hE5, 8'hF0, 8'hC4},
{8'hE6, 8'hE6, 8'hCB},
{8'hEF, 8'hE2, 8'hDA},
{8'hC0, 8'hA7, 8'hA5},
{8'hB7, 8'h9B, 8'h94},
{8'hD2, 8'hC0, 8'hB4},
{8'hFC, 8'hF6, 8'hEF},
{8'hFD, 8'hFB, 8'hF7},
{8'hE7, 8'hE3, 8'hC5},
{8'hE6, 8'hDB, 8'hC4},
{8'hF3, 8'hE2, 8'hD4},
{8'hC5, 8'hAE, 8'h9E},
{8'hE7, 8'hD5, 8'hBD},
{8'hF4, 8'hEB, 8'hD2},
{8'hFA, 8'hF7, 8'hEB},
{8'hF4, 8'hF4, 8'hF2},
{8'hE9, 8'hE8, 8'hD3},
{8'hD4, 8'hD1, 8'hBD},
{8'hA5, 8'hA3, 8'h8E},
{8'h99, 8'h98, 8'h7A},
{8'h93, 8'h93, 8'h6D},
{8'hBB, 8'hBA, 8'h99},
{8'hD5, 8'hD1, 8'hC4},
{8'h26, 8'h21, 8'h28},
{8'h04, 8'h03, 8'h1D},
{8'h06, 8'h02, 8'h19},
{8'h05, 8'h00, 8'h1A},
{8'h00, 8'h01, 8'h30},
{8'h0A, 8'h2F, 8'h78},
{8'h15, 8'h53, 8'hB2},
{8'h14, 8'h55, 8'hB8},
{8'h1B, 8'h55, 8'hB6},
{8'h17, 8'h51, 8'hB7},
{8'h17, 8'h53, 8'hB2},
{8'h1F, 8'h4F, 8'h9B},
{8'h11, 8'h48, 8'h98},
{8'h0C, 8'h45, 8'h9F},
{8'h4D, 8'h57, 8'h84},
{8'hB7, 8'h9F, 8'hA0},
{8'hBE, 8'hC1, 8'hC5},
{8'hB7, 8'hBB, 8'hBB},
{8'h95, 8'h97, 8'h96},
{8'h6E, 8'h6F, 8'h6E},
{8'h75, 8'h73, 8'h74},
{8'h8F, 8'h8B, 8'h8C},
{8'h73, 8'h6E, 8'h70},
{8'h91, 8'h8B, 8'h8D},
{8'hC5, 8'hBD, 8'hC0},
{8'h7C, 8'h76, 8'h8F},
{8'h00, 8'h00, 8'h0B},
{8'h32, 8'h2F, 8'h35},
{8'hCC, 8'hC8, 8'hBD},
{8'hEA, 8'hE6, 8'hCA},
{8'hEE, 8'hE8, 8'hC1},
{8'hDB, 8'hD4, 8'hA6},
{8'hE2, 8'hDB, 8'hAA},
{8'hE3, 8'hDF, 8'hBF},
{8'hEC, 8'hE7, 8'hD5},
{8'hF7, 8'hF1, 8'hED},
{8'hF7, 8'hF2, 8'hEE},
{8'hF9, 8'hF7, 8'hE8},
{8'hF9, 8'hF9, 8'hE4},
{8'hF3, 8'hF5, 8'hE3},
{8'hF6, 8'hF6, 8'hEC},
{8'hEE, 8'hEE, 8'hDC},
{8'hE7, 8'hE6, 8'hCD},
{8'hF2, 8'hEC, 8'hD7},
{8'hE7, 8'hDE, 8'hC4},
{8'hD9, 8'hD2, 8'h8F},
{8'hDC, 8'hD7, 8'h68},
{8'hEB, 8'hE0, 8'h7D},
{8'hFA, 8'hE8, 8'hB5},
{8'hF9, 8'hF3, 8'hCD},
{8'hF7, 8'hF3, 8'hD3},
{8'hF4, 8'hF1, 8'hDC},
{8'hEE, 8'hEC, 8'hDF},
{8'hE3, 8'hE5, 8'hD5},
{8'hD4, 8'hDA, 8'hBD},
{8'hE7, 8'hF2, 8'hC6},
{8'hE0, 8'hF0, 8'hB7},
{8'hE0, 8'hEE, 8'hB4},
{8'hEA, 8'hF6, 8'hC3},
{8'hC1, 8'hCC, 8'hA2},
{8'hB1, 8'hBB, 8'h9A},
{8'hD4, 8'hDD, 8'hC3},
{8'h88, 8'h90, 8'h7A},
{8'h89, 8'h90, 8'h7B},
{8'hB6, 8'hBD, 8'hA9},
{8'hE4, 8'hF3, 8'hD2},
{8'hEA, 8'hFB, 8'hBF},
{8'hD5, 8'hE0, 8'hB8},
{8'h69, 8'h67, 8'h6E},
{8'h14, 8'h06, 8'h09},
{8'h65, 8'h3E, 8'h0F},
{8'h98, 8'h55, 8'h1F},
{8'h60, 8'h0C, 8'h0A},
{8'h50, 8'h3A, 8'h35},
{8'h86, 8'h7B, 8'h78},
{8'h82, 8'h7E, 8'h81},
{8'h7B, 8'h7C, 8'h83},
{8'h7D, 8'h7D, 8'h84},
{8'h7C, 8'h78, 8'h7B},
{8'h8C, 8'h80, 8'h7E},
{8'h88, 8'h77, 8'h70},
{8'h87, 8'h72, 8'h6E},
{8'h85, 8'h70, 8'h6C},
{8'h84, 8'h6E, 8'h6A},
{8'h85, 8'h70, 8'h6B},
{8'h8E, 8'h79, 8'h75},
{8'h87, 8'h72, 8'h6D},
{8'h87, 8'h72, 8'h6D},
{8'h89, 8'h72, 8'h6E},
{8'hA5, 8'h7D, 8'h7C},
{8'hD1, 8'hA4, 8'hA0},
{8'hF5, 8'hC9, 8'hC0},
{8'hF5, 8'hC8, 8'hBA},
{8'hE4, 8'hAE, 8'hA0},
{8'hEC, 8'hB8, 8'hAE},
{8'hB2, 8'h84, 8'h81},
{8'h94, 8'h6C, 8'h6D},
{8'h7F, 8'h7D, 8'h7E},
{8'h7F, 8'h7D, 8'h7E},
{8'h7F, 8'h7D, 8'h7E},
{8'h7F, 8'h7D, 8'h7E},
{8'h80, 8'h7E, 8'h7F},
{8'h7F, 8'h7D, 8'h7E},
{8'h85, 8'h83, 8'h84},
{8'h8D, 8'h8C, 8'h8D},
{8'h92, 8'h92, 8'h95},
{8'h8F, 8'h8E, 8'h94},
{8'h89, 8'h89, 8'h87},
{8'h88, 8'h8B, 8'h76},
{8'hD1, 8'hD9, 8'hAD},
{8'hED, 8'hF6, 8'hBF},
{8'hE9, 8'hF2, 8'hC1},
{8'hE9, 8'hF1, 8'hC8},
{8'hDC, 8'hEB, 8'hBB},
{8'hED, 8'hF1, 8'hD5},
{8'hE7, 8'hDE, 8'hD9},
{8'hE6, 8'hD2, 8'hD9},
{8'hE5, 8'hD3, 8'hD3},
{8'hFC, 8'hF4, 8'hEA},
{8'hF3, 8'hF2, 8'hE6},
{8'hF8, 8'hFA, 8'hEE},
{8'hE2, 8'hDF, 8'hC4},
{8'hEF, 8'hE6, 8'hD4},
{8'hFD, 8'hF0, 8'hE4},
{8'hEE, 8'hDB, 8'hCC},
{8'hDD, 8'hCC, 8'hB2},
{8'hE8, 8'hDF, 8'hC1},
{8'hFC, 8'hF9, 8'hE5},
{8'hEC, 8'hEB, 8'hDE},
{8'hE1, 8'hE2, 8'hBC},
{8'hDA, 8'hD9, 8'hBB},
{8'hA0, 8'h9D, 8'h89},
{8'h92, 8'h90, 8'h79},
{8'hAF, 8'hAF, 8'h8F},
{8'h96, 8'h96, 8'h71},
{8'hDB, 8'hD9, 8'hBC},
{8'h9A, 8'h99, 8'h88},
{8'h01, 8'h03, 8'h18},
{8'h04, 8'h02, 8'h1A},
{8'h09, 8'h02, 8'h18},
{8'h03, 8'h01, 8'h20},
{8'h01, 8'h0B, 8'h41},
{8'h17, 8'h43, 8'h92},
{8'h18, 8'h53, 8'hB0},
{8'h13, 8'h53, 8'hB6},
{8'h10, 8'h52, 8'hB9},
{8'h0E, 8'h56, 8'hB9},
{8'h0F, 8'h57, 8'hB3},
{8'h0C, 8'h58, 8'hBB},
{8'h10, 8'h53, 8'hBA},
{8'h42, 8'h59, 8'h9A},
{8'hCE, 8'hBE, 8'hD2},
{8'hCA, 8'hC0, 8'hC5},
{8'hB6, 8'hB5, 8'hB6},
{8'hA3, 8'hA3, 8'hA3},
{8'hA2, 8'hA1, 8'hA1},
{8'hC2, 8'hC1, 8'hC2},
{8'hC9, 8'hC7, 8'hC8},
{8'hB0, 8'hAD, 8'hAE},
{8'h9C, 8'h97, 8'h98},
{8'hA2, 8'h9D, 8'h9F},
{8'h79, 8'h74, 8'h8D},
{8'h0A, 8'h06, 8'h1F},
{8'h25, 8'h20, 8'h2E},
{8'hD5, 8'hCF, 8'hD0},
{8'hEC, 8'hE6, 8'hDB},
{8'hED, 8'hE6, 8'hD2},
{8'hE2, 8'hDB, 8'hC0},
{8'hDE, 8'hD6, 8'hB8},
{8'hE4, 8'hE0, 8'hC3},
{8'hEF, 8'hEB, 8'hD9},
{8'hED, 8'hE9, 8'hDE},
{8'hF0, 8'hED, 8'hDE},
{8'hE0, 8'hE1, 8'hC4},
{8'hCC, 8'hD0, 8'hA9},
{8'hD6, 8'hDB, 8'hB7},
{8'hE1, 8'hE4, 8'hC8},
{8'hEB, 8'hEA, 8'hD0},
{8'hEA, 8'hE8, 8'hCF},
{8'hEF, 8'hEC, 8'hDA},
{8'hF8, 8'hF3, 8'hDE},
{8'hE8, 8'hE5, 8'hB5},
{8'hE8, 8'hE7, 8'h9E},
{8'hEE, 8'hEA, 8'hAD},
{8'hF5, 8'hEC, 8'hCE},
{8'hF4, 8'hEE, 8'hD7},
{8'hFE, 8'hF9, 8'hE6},
{8'hFA, 8'hF6, 8'hE8},
{8'hE9, 8'hE7, 8'hDB},
{8'hD6, 8'hD8, 8'hC5},
{8'h8F, 8'h95, 8'h75},
{8'hA6, 8'hB0, 8'h83},
{8'hE2, 8'hEF, 8'hB8},
{8'hE8, 8'hF5, 8'hBC},
{8'hDF, 8'hEC, 8'hB6},
{8'hBD, 8'hC9, 8'h9A},
{8'hB7, 8'hC2, 8'h99},
{8'hDB, 8'hE5, 8'hBF},
{8'hA3, 8'hAE, 8'h88},
{8'hBE, 8'hC9, 8'hA1},
{8'hDA, 8'hE5, 8'hBC},
{8'hDF, 8'hF2, 8'hC3},
{8'hE0, 8'hF6, 8'hB1},
{8'hE6, 8'hF7, 8'hC2},
{8'hEE, 8'hED, 8'hE2},
{8'hB8, 8'hA5, 8'h99},
{8'h79, 8'h55, 8'h27},
{8'h96, 8'h57, 8'h20},
{8'h67, 8'h19, 8'h0F},
{8'h68, 8'h58, 8'h54},
{8'h85, 8'h80, 8'h7E},
{8'h7D, 8'h7D, 8'h7F},
{8'h7A, 8'h7D, 8'h83},
{8'h79, 8'h7C, 8'h81},
{8'h83, 8'h82, 8'h85},
{8'h83, 8'h7D, 8'h7A},
{8'h85, 8'h7B, 8'h76},
{8'h7B, 8'h78, 8'h7D},
{8'h80, 8'h7D, 8'h83},
{8'h82, 8'h7F, 8'h84},
{8'h80, 8'h7D, 8'h82},
{8'h81, 8'h7E, 8'h83},
{8'h80, 8'h7D, 8'h83},
{8'h80, 8'h7D, 8'h82},
{8'h82, 8'h7D, 8'h82},
{8'h8F, 8'h78, 8'h76},
{8'h8F, 8'h71, 8'h6C},
{8'h95, 8'h70, 8'h66},
{8'hAE, 8'h84, 8'h74},
{8'hA6, 8'h7B, 8'h6B},
{8'h8D, 8'h64, 8'h56},
{8'h93, 8'h6E, 8'h63},
{8'h8E, 8'h6C, 8'h64},
{8'h7F, 8'h7D, 8'h7E},
{8'h7F, 8'h7D, 8'h7E},
{8'h7E, 8'h7C, 8'h7D},
{8'h7E, 8'h7C, 8'h7D},
{8'h81, 8'h7F, 8'h80},
{8'h7E, 8'h7C, 8'h7D},
{8'h7F, 8'h7D, 8'h7D},
{8'h7C, 8'h7B, 8'h7C},
{8'h7A, 8'h78, 8'h84},
{8'h7C, 8'h7B, 8'h84},
{8'h76, 8'h77, 8'h70},
{8'h8F, 8'h95, 8'h74},
{8'hEA, 8'hF2, 8'hBD},
{8'hEC, 8'hF4, 8'hBC},
{8'hEE, 8'hF4, 8'hCB},
{8'hB0, 8'hB5, 8'h9A},
{8'hB4, 8'hC4, 8'h95},
{8'hEF, 8'hF8, 8'hDC},
{8'hED, 8'hE8, 8'hE6},
{8'hED, 8'hE0, 8'hE7},
{8'hF8, 8'hEC, 8'hEC},
{8'hF4, 8'hEF, 8'hE2},
{8'hFA, 8'hFA, 8'hEB},
{8'hF7, 8'hFA, 8'hEC},
{8'hDB, 8'hDA, 8'hC2},
{8'hED, 8'hE7, 8'hD7},
{8'hFE, 8'hF6, 8'hEF},
{8'hFA, 8'hEE, 8'hE1},
{8'hDA, 8'hCE, 8'hB5},
{8'hDE, 8'hD8, 8'hB8},
{8'hFC, 8'hF9, 8'hDF},
{8'hE8, 8'hE6, 8'hD2},
{8'hEE, 8'hEE, 8'hCA},
{8'hD7, 8'hD5, 8'hBE},
{8'hBC, 8'hB8, 8'hB0},
{8'hCA, 8'hC6, 8'hBE},
{8'hD8, 8'hD5, 8'hC2},
{8'h8F, 8'h8E, 8'h6F},
{8'hB2, 8'hB1, 8'h91},
{8'hDC, 8'hDC, 8'hC4},
{8'h3D, 8'h46, 8'h5C},
{8'h00, 8'h00, 8'h11},
{8'h0B, 8'h06, 8'h17},
{8'h08, 8'h02, 8'h16},
{8'h02, 8'h01, 8'h25},
{8'h08, 8'h1A, 8'h56},
{8'h18, 8'h4A, 8'h9D},
{8'h15, 8'h55, 8'hB7},
{8'h0E, 8'h56, 8'hC0},
{8'h0E, 8'h57, 8'hBA},
{8'h13, 8'h58, 8'hB2},
{8'h19, 8'h54, 8'hAD},
{8'h1E, 8'h47, 8'h9C},
{8'h25, 8'h34, 8'h75},
{8'h66, 8'h61, 8'h84},
{8'h98, 8'h8D, 8'h9B},
{8'hD2, 8'hCF, 8'hD0},
{8'hF5, 8'hF4, 8'hF5},
{8'hF7, 8'hF6, 8'hF7},
{8'hFF, 8'hFF, 8'hFF},
{8'hFF, 8'hFF, 8'hFF},
{8'hFF, 8'hFF, 8'hFF},
{8'hFD, 8'hFC, 8'hFD},
{8'hD3, 8'hD0, 8'hD3},
{8'h87, 8'h83, 8'h97},
{8'h1C, 8'h19, 8'h2A},
{8'h38, 8'h33, 8'h3E},
{8'hD0, 8'hCB, 8'hCC},
{8'hF3, 8'hEE, 8'hE6},
{8'hEE, 8'hE9, 8'hD9},
{8'hE8, 8'hE3, 8'hCC},
{8'hE3, 8'hDD, 8'hC3},
{8'hEB, 8'hE9, 8'hD0},
{8'hE9, 8'hE6, 8'hD5},
{8'hF3, 8'hF1, 8'hE4},
{8'hDC, 8'hDC, 8'hC4},
{8'hBE, 8'hC2, 8'h9A},
{8'hBB, 8'hC2, 8'h8F},
{8'hE1, 8'hE8, 8'hB8},
{8'hD5, 8'hDC, 8'hB3},
{8'hDB, 8'hDA, 8'hBB},
{8'hEA, 8'hE8, 8'hD2},
{8'hF0, 8'hEC, 8'hDF},
{8'hF8, 8'hF5, 8'hE3},
{8'hEE, 8'hEE, 8'hD1},
{8'hEE, 8'hEF, 8'hCC},
{8'hF6, 8'hF5, 8'hDB},
{8'hFD, 8'hFA, 8'hED},
{8'hF8, 8'hF5, 8'hEA},
{8'hF9, 8'hF5, 8'hEA},
{8'hFD, 8'hFD, 8'hF1},
{8'hFD, 8'hFC, 8'hEF},
{8'hEA, 8'hEC, 8'hD5},
{8'h8E, 8'h93, 8'h70},
{8'h87, 8'h8F, 8'h62},
{8'hDE, 8'hE8, 8'hB4},
{8'hE8, 8'hF5, 8'hBE},
{8'hD5, 8'hE2, 8'hAD},
{8'hA7, 8'hB3, 8'h82},
{8'hD4, 8'hE0, 8'hB2},
{8'hE5, 8'hF1, 8'hC3},
{8'hE4, 8'hF1, 8'hBF},
{8'hE9, 8'hF6, 8'hC1},
{8'hE7, 8'hF2, 8'hBD},
{8'hE3, 8'hF2, 8'hB8},
{8'hE5, 8'hF9, 8'hB2},
{8'hDF, 8'hF1, 8'hB7},
{8'hE5, 8'hF0, 8'hCF},
{8'hF1, 8'hF2, 8'hCA},
{8'hEE, 8'hE5, 8'hA0},
{8'hB3, 8'h99, 8'h5D},
{8'h5E, 8'h38, 8'h21},
{8'h74, 8'h6C, 8'h68},
{8'h81, 8'h7F, 8'h7E},
{8'h7D, 8'h7E, 8'h7F},
{8'h7B, 8'h80, 8'h83},
{8'h7B, 8'h7F, 8'h83},
{8'h7F, 8'h80, 8'h81},
{8'h81, 8'h7E, 8'h7C},
{8'h82, 8'h7E, 8'h7A},
{8'h7D, 8'h7E, 8'h83},
{8'h7D, 8'h7F, 8'h84},
{8'h7D, 8'h7E, 8'h84},
{8'h7C, 8'h7E, 8'h83},
{8'h7B, 8'h7D, 8'h82},
{8'h7C, 8'h7D, 8'h83},
{8'h7D, 8'h7F, 8'h84},
{8'h7B, 8'h7D, 8'h82},
{8'h77, 8'h7E, 8'h7F},
{8'h79, 8'h7D, 8'h7A},
{8'h80, 8'h7F, 8'h77},
{8'h80, 8'h7A, 8'h6F},
{8'h7D, 8'h74, 8'h67},
{8'h85, 8'h7B, 8'h6E},
{8'h7B, 8'h73, 8'h67},
{8'h83, 8'h7D, 8'h72},
{8'h7E, 8'h7C, 8'h7D},
{8'h7E, 8'h7C, 8'h7D},
{8'h7E, 8'h7C, 8'h7D},
{8'h7F, 8'h7D, 8'h7E},
{8'h7F, 8'h7D, 8'h7E},
{8'h7D, 8'h7B, 8'h7C},
{8'h7E, 8'h7C, 8'h7C},
{8'h82, 8'h80, 8'h82},
{8'h7C, 8'h79, 8'h86},
{8'h8C, 8'h89, 8'h92},
{8'h8C, 8'h8D, 8'h86},
{8'hA8, 8'hAD, 8'h8D},
{8'hEC, 8'hF4, 8'hC1},
{8'hF0, 8'hF7, 8'hC6},
{8'hC4, 8'hC8, 8'hAB},
{8'h75, 8'h78, 8'h6B},
{8'h98, 8'hA8, 8'h7F},
{8'hE2, 8'hEB, 8'hD0},
{8'hE5, 8'hE4, 8'hDD},
{8'hE9, 8'hE3, 8'hE0},
{8'hF4, 8'hEE, 8'hE3},
{8'hE6, 8'hE3, 8'hCF},
{8'hE4, 8'hE6, 8'hD2},
{8'hF2, 8'hF5, 8'hE6},
{8'hCC, 8'hCD, 8'hB6},
{8'hEA, 8'hE7, 8'hDA},
{8'hFC, 8'hF6, 8'hF2},
{8'hFE, 8'hF7, 8'hF0},
{8'hF4, 8'hEF, 8'hDB},
{8'hD2, 8'hCD, 8'hB1},
{8'hE4, 8'hE0, 8'hC7},
{8'hE9, 8'hE4, 8'hD2},
{8'hF0, 8'hEE, 8'hDA},
{8'hF9, 8'hF5, 8'hEE},
{8'hFF, 8'hF8, 8'hFE},
{8'hFE, 8'hF8, 8'hFD},
{8'hF8, 8'hF4, 8'hEA},
{8'hBF, 8'hBD, 8'hA7},
{8'hA3, 8'hA0, 8'h87},
{8'hBF, 8'hBE, 8'hAA},
{8'hBE, 8'hC6, 8'hCD},
{8'h0E, 8'h11, 8'h1F},
{8'h04, 8'h04, 8'h10},
{8'h06, 8'h01, 8'h0E},
{8'h07, 8'h01, 8'h19},
{8'h00, 8'h00, 8'h2B},
{8'h12, 8'h32, 8'h79},
{8'h1E, 8'h58, 8'hB3},
{8'h0E, 8'h53, 8'hB8},
{8'h19, 8'h58, 8'hB0},
{8'h19, 8'h50, 8'h9C},
{8'h2E, 8'h4E, 8'h90},
{8'h3C, 8'h42, 8'h7A},
{8'h1D, 8'h24, 8'h5F},
{8'h7C, 8'h86, 8'hB4},
{8'hF1, 8'hEA, 8'hFA},
{8'hFF, 8'hFF, 8'hFF},
{8'hFD, 8'hFC, 8'hFD},
{8'hE8, 8'hE5, 8'hE6},
{8'hFD, 8'hFC, 8'hFD},
{8'hFE, 8'hFD, 8'hFE},
{8'hFB, 8'hFA, 8'hFB},
{8'hFB, 8'hFB, 8'hFB},
{8'hFB, 8'hFA, 8'hFB},
{8'hCD, 8'hCA, 8'hD3},
{8'h50, 8'h4D, 8'h55},
{8'h68, 8'h64, 8'h69},
{8'hBF, 8'hBB, 8'hB9},
{8'hF2, 8'hEF, 8'hE5},
{8'hEB, 8'hEA, 8'hD7},
{8'hF0, 8'hEE, 8'hD3},
{8'hDF, 8'hDE, 8'hBF},
{8'hEF, 8'hEE, 8'hD9},
{8'hEA, 8'hE8, 8'hDA},
{8'hFB, 8'hFA, 8'hEC},
{8'hD6, 8'hD8, 8'hBE},
{8'hB8, 8'hBF, 8'h91},
{8'hDA, 8'hE4, 8'hAC},
{8'hED, 8'hF6, 8'hC3},
{8'hC7, 8'hD0, 8'hA4},
{8'hBE, 8'hBF, 8'h9D},
{8'hDA, 8'hD8, 8'hC6},
{8'hEC, 8'hE9, 8'hDF},
{8'hF9, 8'hF9, 8'hE7},
{8'hF6, 8'hF5, 8'hE3},
{8'hF4, 8'hF1, 8'hEA},
{8'hF9, 8'hF7, 8'hF4},
{8'hFF, 8'hFF, 8'hF5},
{8'hFD, 8'hFC, 8'hF5},
{8'hFB, 8'hFA, 8'hF0},
{8'hF9, 8'hF8, 8'hEA},
{8'hF7, 8'hF8, 8'hE2},
{8'hF4, 8'hF7, 8'hD8},
{8'hD7, 8'hDB, 8'hB5},
{8'hD3, 8'hD9, 8'hAE},
{8'hD5, 8'hDD, 8'hAD},
{8'hC7, 8'hD4, 8'h9F},
{8'hCA, 8'hD6, 8'hA3},
{8'hD2, 8'hDE, 8'hAF},
{8'hD4, 8'hE0, 8'hB2},
{8'hD4, 8'hE0, 8'hB0},
{8'hDE, 8'hEB, 8'hB7},
{8'hE5, 8'hF3, 8'hBA},
{8'hE6, 8'hF4, 8'hB8},
{8'hEA, 8'hF1, 8'hB5},
{8'hE7, 8'hF2, 8'hB2},
{8'hE3, 8'hF4, 8'hBA},
{8'hDF, 8'hF4, 8'hC2},
{8'hDB, 8'hF3, 8'hB8},
{8'hE1, 8'hF8, 8'hAF},
{8'hEE, 8'hFC, 8'hC0},
{8'hA5, 8'hAD, 8'h8A},
{8'h7E, 8'h7D, 8'h7A},
{8'h7F, 8'h7F, 8'h80},
{8'h7E, 8'h7F, 8'h81},
{8'h7D, 8'h7E, 8'h81},
{8'h7D, 8'h7E, 8'h81},
{8'h7D, 8'h7E, 8'h80},
{8'h7F, 8'h7E, 8'h7F},
{8'h7F, 8'h7D, 8'h7D},
{8'h80, 8'h7D, 8'h7E},
{8'h80, 8'h7D, 8'h7E},
{8'h80, 8'h7D, 8'h7E},
{8'h80, 8'h7D, 8'h7E},
{8'h80, 8'h7D, 8'h7E},
{8'h80, 8'h7D, 8'h7E},
{8'h80, 8'h7C, 8'h7E},
{8'h7F, 8'h7D, 8'h7F},
{8'h79, 8'h7E, 8'h89},
{8'h7A, 8'h7E, 8'h89},
{8'h7D, 8'h7D, 8'h85},
{8'h7F, 8'h7D, 8'h83},
{8'h81, 8'h7D, 8'h80},
{8'h82, 8'h7C, 8'h7F},
{8'h83, 8'h7D, 8'h80},
{8'h81, 8'h7C, 8'h7F},
{8'h7F, 8'h7D, 8'h7E},
{8'h7D, 8'h7B, 8'h7C},
{8'h7F, 8'h7D, 8'h7E},
{8'h84, 8'h82, 8'h83},
{8'h7E, 8'h7C, 8'h7D},
{8'h7C, 8'h7A, 8'h7B},
{8'h7F, 8'h7D, 8'h7E},
{8'h77, 8'h75, 8'h76},
{8'hB3, 8'hB2, 8'hB6},
{8'hEA, 8'hE9, 8'hED},
{8'hC0, 8'hC1, 8'hBC},
{8'hCE, 8'hD1, 8'hBA},
{8'hF3, 8'hF9, 8'hD4},
{8'hCA, 8'hD0, 8'hAC},
{8'h80, 8'h82, 8'h71},
{8'h79, 8'h79, 8'h77},
{8'h8C, 8'h97, 8'h79},
{8'hDA, 8'hDF, 8'hC9},
{8'hD8, 8'hD8, 8'hC8},
{8'hDF, 8'hDC, 8'hC9},
{8'hE8, 8'hE6, 8'hC9},
{8'hE6, 8'hE5, 8'hC6},
{8'hEB, 8'hEA, 8'hD7},
{8'hF2, 8'hF2, 8'hE8},
{8'hC5, 8'hC8, 8'hB1},
{8'hE1, 8'hE2, 8'hD6},
{8'hFF, 8'hFD, 8'hFC},
{8'hFA, 8'hF7, 8'hF5},
{8'hFF, 8'hFE, 8'hF2},
{8'hEA, 8'hE6, 8'hD2},
{8'hD0, 8'hCA, 8'hB9},
{8'hF4, 8'hEC, 8'hE3},
{8'hFB, 8'hF6, 8'hF0},
{8'hF8, 8'hF2, 8'hF5},
{8'hFB, 8'hF4, 8'hFD},
{8'hFC, 8'hF7, 8'hF8},
{8'hF0, 8'hEE, 8'hDF},
{8'hD0, 8'hCE, 8'hB5},
{8'hC7, 8'hC5, 8'hAF},
{8'hDA, 8'hD7, 8'hC8},
{8'hF5, 8'hF5, 8'hF4},
{8'h7C, 8'h80, 8'h87},
{8'h00, 8'h01, 8'h0B},
{8'h04, 8'h03, 8'h12},
{8'h07, 8'h01, 8'h11},
{8'h05, 8'h01, 8'h22},
{8'h07, 8'h14, 8'h4D},
{8'h26, 8'h52, 8'hA0},
{8'h24, 8'h52, 8'hA5},
{8'h11, 8'h3A, 8'h83},
{8'h06, 8'h34, 8'h7A},
{8'h46, 8'h61, 8'h9C},
{8'h88, 8'h86, 8'hB3},
{8'h32, 8'h42, 8'h7C},
{8'h65, 8'h7E, 8'hB0},
{8'hFF, 8'hFC, 8'hFF},
{8'hFF, 8'hFF, 8'hFF},
{8'hFA, 8'hF5, 8'hF7},
{8'hE8, 8'hE4, 8'hE5},
{8'hFF, 8'hFF, 8'hFF},
{8'hFF, 8'hFF, 8'hFF},
{8'hFF, 8'hFF, 8'hFF},
{8'hFF, 8'hFF, 8'hFF},
{8'hFC, 8'hFC, 8'hFC},
{8'hD4, 8'hCF, 8'hDA},
{8'h5D, 8'h58, 8'h63},
{8'h37, 8'h33, 8'h3A},
{8'h7A, 8'h78, 8'h7A},
{8'hF9, 8'hF8, 8'hF2},
{8'hED, 8'hEE, 8'hDC},
{8'hD6, 8'hD9, 8'hBC},
{8'hE4, 8'hE7, 8'hC6},
{8'hE0, 8'hDE, 8'hCF},
{8'hF1, 8'hF0, 8'hE6},
{8'hF3, 8'hF3, 8'hE7},
{8'hEB, 8'hEE, 8'hD5},
{8'hD3, 8'hDB, 8'hAE},
{8'hEA, 8'hF4, 8'hBF},
{8'hE3, 8'hEC, 8'hBF},
{8'hA7, 8'hB0, 8'h8C},
{8'hB7, 8'hB9, 8'h97},
{8'hDD, 8'hDC, 8'hCF},
{8'hF3, 8'hF1, 8'hE8},
{8'hF6, 8'hF5, 8'hE0},
{8'hFB, 8'hF8, 8'hEA},
{8'hFC, 8'hF4, 8'hFD},
{8'hFD, 8'hF5, 8'hFB},
{8'hFE, 8'hFA, 8'hE9},
{8'hF9, 8'hF9, 8'hEE},
{8'hF6, 8'hF6, 8'hE8},
{8'hF2, 8'hF5, 8'hDD},
{8'hF9, 8'hFC, 8'hDC},
{8'hE1, 8'hE6, 8'hBF},
{8'hDC, 8'hE0, 8'hB6},
{8'hD3, 8'hD7, 8'hAE},
{8'hD3, 8'hD7, 8'hAD},
{8'hDD, 8'hE8, 8'hB8},
{8'hE5, 8'hF1, 8'hC2},
{8'hE7, 8'hF2, 8'hC6},
{8'hE2, 8'hED, 8'hC3},
{8'hE0, 8'hEC, 8'hC1},
{8'hE2, 8'hEE, 8'hC0},
{8'hE3, 8'hF0, 8'hBD},
{8'hE4, 8'hF0, 8'hB9},
{8'hE9, 8'hF1, 8'hB6},
{8'hE7, 8'hF2, 8'hB9},
{8'hE3, 8'hF3, 8'hBE},
{8'hDE, 8'hF5, 8'hBB},
{8'hDC, 8'hF8, 8'hB8},
{8'hDA, 8'hF8, 8'hB7},
{8'hE1, 8'hFC, 8'hC9},
{8'hD6, 8'hEC, 8'hCC},
{8'h85, 8'h84, 8'h86},
{8'h7F, 8'h7D, 8'h81},
{8'h80, 8'h7D, 8'h80},
{8'h80, 8'h7D, 8'h80},
{8'h80, 8'h7D, 8'h80},
{8'h80, 8'h7D, 8'h80},
{8'hFF, 8'hD7, 8'h00},
{8'h7F, 8'h7D, 8'h81},
{8'h82, 8'h7C, 8'h7C},
{8'h82, 8'h7C, 8'h7C},
{8'h82, 8'h7C, 8'h7C},
{8'h82, 8'h7C, 8'h7C},
{8'h82, 8'h7C, 8'h7C},
{8'h82, 8'h7C, 8'h7C},
{8'h82, 8'h7C, 8'h7C},
{8'h83, 8'h7C, 8'h7D},
{8'h86, 8'h78, 8'h87},
{8'h87, 8'h78, 8'h87},
{8'h87, 8'h78, 8'h87},
{8'h87, 8'h78, 8'h87},
{8'h87, 8'h77, 8'h87},
{8'h87, 8'h77, 8'h86},
{8'h88, 8'h78, 8'h85},
{8'h88, 8'h78, 8'h85},
{8'h89, 8'h87, 8'h89},
{8'h7F, 8'h7D, 8'h7E},
{8'h7B, 8'h79, 8'h7B},
{8'h81, 8'h7F, 8'h80},
{8'h80, 8'h7E, 8'h7F},
{8'h7C, 8'h7A, 8'h7B},
{8'h90, 8'h8E, 8'h8F},
{8'hA5, 8'hA3, 8'hA3},
{8'hDC, 8'hDE, 8'hD7},
{8'hF0, 8'hF0, 8'hEE},
{8'hCF, 8'hCF, 8'hCD},
{8'hE6, 8'hE8, 8'hDC},
{8'hCF, 8'hD3, 8'hBB},
{8'h8E, 8'h91, 8'h7B},
{8'h87, 8'h89, 8'h82},
{8'hA5, 8'hA4, 8'hAB},
{8'hE9, 8'hEC, 8'hDA},
{8'hEA, 8'hEC, 8'hD8},
{8'hEC, 8'hED, 8'hD4},
{8'hD7, 8'hD8, 8'hB2},
{8'hBC, 8'hBC, 8'h8B},
{8'hCD, 8'hCB, 8'hA2},
{8'hF3, 8'hF0, 8'hDC},
{8'hE9, 8'hE5, 8'hE2},
{8'hC9, 8'hCD, 8'hB5},
{8'hD6, 8'hD8, 8'hCB},
{8'hF9, 8'hFA, 8'hFC},
{8'hF5, 8'hF5, 8'hFA},
{8'hF7, 8'hF5, 8'hF1},
{8'hF6, 8'hF2, 8'hE7},
{8'hE4, 8'hDD, 8'hD6},
{8'hF8, 8'hEF, 8'hEE},
{8'hFB, 8'hF4, 8'hF4},
{8'hFA, 8'hF4, 8'hF7},
{8'hFB, 8'hF5, 8'hF5},
{8'hF7, 8'hF5, 8'hE6},
{8'hC8, 8'hC7, 8'hA7},
{8'hC5, 8'hC6, 8'hA0},
{8'hDC, 8'hDA, 8'hBF},
{8'hF3, 8'hEF, 8'hDE},
{8'hF8, 8'hEE, 8'hE2},
{8'hE6, 8'hE9, 8'hE9},
{8'h29, 8'h33, 8'h41},
{8'h01, 8'h04, 8'h15},
{8'h08, 8'h02, 8'h12},
{8'h09, 8'h03, 8'h1E},
{8'h02, 8'h09, 8'h3A},
{8'h11, 8'h2F, 8'h72},
{8'h0B, 8'h17, 8'h51},
{8'h06, 8'h17, 8'h4F},
{8'h16, 8'h4F, 8'h9A},
{8'h2B, 8'h5A, 8'hA0},
{8'h52, 8'h62, 8'h97},
{8'h15, 8'h34, 8'h78},
{8'h36, 8'h57, 8'h8A},
{8'hB6, 8'hAB, 8'hA2},
{8'hB2, 8'hAC, 8'hAB},
{8'h9A, 8'h92, 8'h95},
{8'h96, 8'h91, 8'h92},
{8'hA2, 8'h9F, 8'h9F},
{8'hB2, 8'hB1, 8'hB2},
{8'hAB, 8'hAC, 8'hAB},
{8'h86, 8'h89, 8'h87},
{8'h79, 8'h7B, 8'h7B},
{8'h8F, 8'h88, 8'h99},
{8'h89, 8'h7F, 8'h97},
{8'h16, 8'h11, 8'h25},
{8'h21, 8'h1F, 8'h2D},
{8'hE3, 8'hE1, 8'hE6},
{8'hF1, 8'hF2, 8'hE8},
{8'hB4, 8'hB7, 8'h9F},
{8'hBC, 8'hC1, 8'hA3},
{8'hAE, 8'hAE, 8'hA2},
{8'hD6, 8'hD6, 8'hD1},
{8'hF0, 8'hF0, 8'hE9},
{8'hED, 8'hF1, 8'hDB},
{8'hE3, 8'hEA, 8'hC3},
{8'hDC, 8'hE5, 8'hB7},
{8'hBD, 8'hC8, 8'hA3},
{8'h9B, 8'hA3, 8'h89},
{8'hDC, 8'hE1, 8'hC0},
{8'hE6, 8'hE6, 8'hDE},
{8'hF3, 8'hF1, 8'hEB},
{8'hF9, 8'hF7, 8'hDE},
{8'hFF, 8'hF9, 8'hEC},
{8'hFF, 8'hF2, 8'hFF},
{8'hFD, 8'hEF, 8'hF6},
{8'hF5, 8'hEE, 8'hD1},
{8'hF6, 8'hF8, 8'hE6},
{8'hEF, 8'hF3, 8'hDE},
{8'hD1, 8'hD5, 8'hB6},
{8'hC1, 8'hC5, 8'h9D},
{8'hD0, 8'hD4, 8'hA7},
{8'hD0, 8'hD3, 8'hA6},
{8'hDA, 8'hDC, 8'hB3},
{8'hE9, 8'hEB, 8'hC4},
{8'hE0, 8'hEC, 8'hBC},
{8'hDF, 8'hEB, 8'hBD},
{8'hDC, 8'hE8, 8'hBE},
{8'hDB, 8'hE6, 8'hC0},
{8'hDE, 8'hE9, 8'hC3},
{8'hDC, 8'hE7, 8'hBF},
{8'hDF, 8'hEA, 8'hBF},
{8'hE4, 8'hF0, 8'hC0},
{8'hE4, 8'hF4, 8'hB8},
{8'hE3, 8'hF2, 8'hC1},
{8'hE2, 8'hF2, 8'hC4},
{8'hE1, 8'hF4, 8'hBA},
{8'hE0, 8'hF1, 8'hB1},
{8'hE0, 8'hED, 8'hBA},
{8'hD7, 8'hDE, 8'hBF},
{8'hAE, 8'hB1, 8'hA0},
{8'h84, 8'h81, 8'h87},
{8'h81, 8'h7C, 8'h82},
{8'h83, 8'h7C, 8'h81},
{8'h83, 8'h7B, 8'h80},
{8'h83, 8'h7B, 8'h80},
{8'h83, 8'h7B, 8'h80},
{8'h81, 8'h7C, 8'h82},
{8'h80, 8'h7C, 8'h83},
{8'h80, 8'h7C, 8'h81},
{8'h80, 8'h7C, 8'h81},
{8'h80, 8'h7C, 8'h81},
{8'h80, 8'h7C, 8'h81},
{8'h80, 8'h7C, 8'h81},
{8'h80, 8'h7C, 8'h81},
{8'h80, 8'h7C, 8'h81},
{8'h81, 8'h7C, 8'h81},
{8'h87, 8'h7A, 8'h7A},
{8'h86, 8'h7A, 8'h7B},
{8'h84, 8'h7B, 8'h7F},
{8'h82, 8'h7B, 8'h82},
{8'h80, 8'h7C, 8'h84},
{8'h80, 8'h7C, 8'h84},
{8'h80, 8'h7C, 8'h83},
{8'h80, 8'h7C, 8'h83},
{8'h90, 8'h8F, 8'h89},
{8'h87, 8'h86, 8'h82},
{8'h78, 8'h76, 8'h76},
{8'h7E, 8'h7C, 8'h7F},
{8'h82, 8'h80, 8'h83},
{8'h7C, 8'h7A, 8'h7D},
{8'hAF, 8'hAD, 8'hAE},
{8'hEB, 8'hEA, 8'hE9},
{8'hD0, 8'hD1, 8'hCC},
{8'hEF, 8'hEF, 8'hEE},
{8'hF6, 8'hF6, 8'hF5},
{8'hFA, 8'hFB, 8'hF4},
{8'hF2, 8'hF3, 8'hE5},
{8'hEE, 8'hEE, 8'hE1},
{8'hE7, 8'hE5, 8'hE2},
{8'hF5, 8'hF2, 8'hF6},
{8'hFA, 8'hF9, 8'hF1},
{8'hF5, 8'hF4, 8'hE7},
{8'hE8, 8'hE6, 8'hCE},
{8'hEF, 8'hEE, 8'hC6},
{8'hE6, 8'hE4, 8'hB5},
{8'hCB, 8'hC8, 8'hA0},
{8'hD7, 8'hD3, 8'hBE},
{8'hEC, 8'hE7, 8'hE2},
{8'hE2, 8'hE6, 8'hD2},
{8'hDD, 8'hE0, 8'hD6},
{8'hEF, 8'hF0, 8'hED},
{8'hF3, 8'hF3, 8'hED},
{8'hF9, 8'hF7, 8'hE8},
{8'hF7, 8'hF2, 8'hE2},
{8'hF1, 8'hE7, 8'hE0},
{8'hF8, 8'hEB, 8'hEE},
{8'hF3, 8'hEF, 8'hEA},
{8'hF3, 8'hEF, 8'hEA},
{8'hFD, 8'hFB, 8'hF2},
{8'hC9, 8'hC8, 8'hB4},
{8'hAF, 8'hB0, 8'h91},
{8'hB7, 8'hB8, 8'h95},
{8'hD1, 8'hD2, 8'hB5},
{8'hF5, 8'hF3, 8'hDC},
{8'hFD, 8'hF5, 8'hE4},
{8'hFC, 8'hFF, 8'hFC},
{8'hAB, 8'hB4, 8'hC2},
{8'h06, 8'h06, 8'h1B},
{8'h08, 8'h02, 8'h14},
{8'h08, 8'h01, 8'h16},
{8'h0E, 8'h15, 8'h38},
{8'h00, 8'h0B, 8'h3A},
{8'h06, 8'h0C, 8'h3D},
{8'h21, 8'h3F, 8'h80},
{8'h19, 8'h53, 8'hA7},
{8'h11, 8'h55, 8'hB6},
{8'h1C, 8'h4F, 8'hA3},
{8'h0A, 8'h3C, 8'h8A},
{8'h15, 8'h45, 8'h7F},
{8'hBE, 8'hC0, 8'hBD},
{8'hCA, 8'hC0, 8'hC4},
{8'h86, 8'h7D, 8'h86},
{8'h65, 8'h5F, 8'h65},
{8'h6C, 8'h6A, 8'h6D},
{8'hA2, 8'hA2, 8'hA2},
{8'hC3, 8'hC5, 8'hC5},
{8'hAE, 8'hB0, 8'hAE},
{8'h9D, 8'h9F, 8'h9F},
{8'h9E, 8'h9B, 8'hAA},
{8'h93, 8'h8E, 8'hA2},
{8'h2A, 8'h23, 8'h3F},
{8'h00, 8'h00, 8'h07},
{8'h8F, 8'h8B, 8'h9B},
{8'hFD, 8'hFC, 8'hF7},
{8'hEA, 8'hEB, 8'hE2},
{8'hB8, 8'hBC, 8'hA9},
{8'h91, 8'h91, 8'h86},
{8'h9C, 8'h9D, 8'h8F},
{8'hD4, 8'hD7, 8'hC0},
{8'hEF, 8'hF4, 8'hD2},
{8'hE4, 8'hEC, 8'hC4},
{8'hC0, 8'hC8, 8'hA2},
{8'hD0, 8'hD7, 8'hBA},
{8'hB7, 8'hBD, 8'hA6},
{8'hD6, 8'hDA, 8'hC4},
{8'hE8, 8'hE9, 8'hDF},
{8'hFA, 8'hFA, 8'hEC},
{8'hE0, 8'hDF, 8'hC6},
{8'hEF, 8'hEA, 8'hDC},
{8'hFD, 8'hF2, 8'hF6},
{8'hF5, 8'hEA, 8'hE5},
{8'hEC, 8'hE6, 8'hC4},
{8'hF1, 8'hF2, 8'hE1},
{8'hB2, 8'hB4, 8'h9D},
{8'hBE, 8'hC4, 8'h9E},
{8'hC8, 8'hCF, 8'h9F},
{8'hD0, 8'hD6, 8'hA5},
{8'hE0, 8'hE5, 8'hBD},
{8'hF4, 8'hF7, 8'hDC},
{8'hF4, 8'hF5, 8'hE1},
{8'hF1, 8'hF8, 8'hDC},
{8'hEC, 8'hF2, 8'hD7},
{8'hE8, 8'hEE, 8'hD3},
{8'hE7, 8'hEC, 8'hD3},
{8'hED, 8'hF4, 8'hDA},
{8'hE5, 8'hEC, 8'hD1},
{8'hDD, 8'hE3, 8'hC7},
{8'hE1, 8'hEA, 8'hC9},
{8'hE0, 8'hF5, 8'hB9},
{8'hE0, 8'hF4, 8'hBE},
{8'hE2, 8'hF2, 8'hC1},
{8'hE4, 8'hF3, 8'hBB},
{8'hEB, 8'hF5, 8'hC0},
{8'hD4, 8'hD9, 8'hB4},
{8'h84, 8'h82, 8'h70},
{8'h7C, 8'h76, 8'h6F},
{8'h81, 8'h7D, 8'h82},
{8'h81, 8'h7D, 8'h82},
{8'h82, 8'h7C, 8'h81},
{8'h83, 8'h7B, 8'h7F},
{8'h83, 8'h7B, 8'h7F},
{8'h82, 8'h7C, 8'h80},
{8'h80, 8'h7C, 8'h81},
{8'h80, 8'h7C, 8'h82},
{8'h7E, 8'h7D, 8'h83},
{8'h7E, 8'h7D, 8'h83},
{8'h7E, 8'h7D, 8'h83},
{8'h7E, 8'h7D, 8'h83},
{8'h7E, 8'h7D, 8'h83},
{8'h7E, 8'h7D, 8'h83},
{8'h7E, 8'h7D, 8'h83},
{8'h7E, 8'h7D, 8'h82},
{8'h81, 8'h7E, 8'h79},
{8'h7F, 8'h7F, 8'h79},
{8'h7D, 8'h7F, 8'h7C},
{8'h7C, 8'h7F, 8'h7E},
{8'h7A, 8'h7F, 8'h80},
{8'h7A, 8'h80, 8'h81},
{8'h7A, 8'h80, 8'h80},
{8'h7A, 8'h80, 8'h80},
{8'h7A, 8'h7A, 8'h72},
{8'h9A, 8'h9A, 8'h92},
{8'h8A, 8'h89, 8'h82},
{8'h79, 8'h78, 8'h72},
{8'h7C, 8'h7B, 8'h77},
{8'h75, 8'h74, 8'h73},
{8'hB1, 8'hAF, 8'hB0},
{8'hE9, 8'hE7, 8'hEA},
{8'hE9, 8'hE8, 8'hEE},
{8'hF1, 8'hF1, 8'hF4},
{8'hFB, 8'hFB, 8'hF7},
{8'hFF, 8'hFF, 8'hF7},
{8'hFF, 8'hFE, 8'hF4},
{8'hFF, 8'hFD, 8'hF4},
{8'hFF, 8'hFB, 8'hF5},
{8'hFC, 8'hF7, 8'hF2},
{8'hFB, 8'hF7, 8'hF1},
{8'hD6, 8'hD2, 8'hC5},
{8'hC3, 8'hBE, 8'hA6},
{8'hEA, 8'hE4, 8'hC5},
{8'hEC, 8'hE6, 8'hC9},
{8'hED, 8'hE9, 8'hD0},
{8'hEC, 8'hE8, 8'hD9},
{8'hF6, 8'hF4, 8'hEB},
{8'hF8, 8'hFB, 8'hF4},
{8'hF4, 8'hF6, 8'hF1},
{8'hEA, 8'hEB, 8'hDF},
{8'hF2, 8'hF1, 8'hD5},
{8'hF2, 8'hF0, 8'hC3},
{8'hF9, 8'hF4, 8'hC7},
{8'hF4, 8'hEA, 8'hCC},
{8'hFA, 8'hEE, 8'hDF},
{8'hF5, 8'hF4, 8'hE6},
{8'hF3, 8'hF3, 8'hE6},
{8'hF4, 8'hF4, 8'hE9},
{8'hEA, 8'hEA, 8'hE1},
{8'hCD, 8'hCD, 8'hC2},
{8'hA1, 8'hA3, 8'h93},
{8'hC6, 8'hC8, 8'hB1},
{8'hEF, 8'hF1, 8'hD6},
{8'hF7, 8'hF7, 8'hE8},
{8'hED, 8'hEF, 8'hED},
{8'hF3, 8'hF5, 8'hFF},
{8'h67, 8'h65, 8'h78},
{8'h05, 8'h00, 8'h0F},
{8'h09, 8'h01, 8'h15},
{8'h05, 8'h06, 8'h1F},
{8'h00, 8'h03, 8'h21},
{8'h15, 8'h33, 8'h75},
{8'h1F, 8'h56, 8'hB4},
{8'h20, 8'h4F, 8'hAC},
{8'h0E, 8'h56, 8'hCA},
{8'h0E, 8'h56, 8'hC4},
{8'h20, 8'h4E, 8'h98},
{8'h12, 8'h45, 8'h83},
{8'h81, 8'h9B, 8'hB9},
{8'h9B, 8'h8C, 8'h9D},
{8'hA1, 8'h94, 8'hA4},
{8'hD4, 8'hCE, 8'hDA},
{8'hFF, 8'hFF, 8'hFF},
{8'hFF, 8'hFF, 8'hFF},
{8'hFF, 8'hFF, 8'hFF},
{8'hFF, 8'hFF, 8'hFF},
{8'hFF, 8'hFF, 8'hFF},
{8'hFA, 8'hFD, 8'hFC},
{8'hD5, 8'hD6, 8'hD9},
{8'h5E, 8'h5B, 8'h6E},
{8'h2A, 8'h27, 8'h2E},
{8'h49, 8'h42, 8'h56},
{8'hE8, 8'hE5, 8'hE4},
{8'hFB, 8'hF9, 8'hF9},
{8'hF4, 8'hF5, 8'hED},
{8'hAE, 8'hB0, 8'hA6},
{8'h9A, 8'h9E, 8'h84},
{8'hC6, 8'hCD, 8'hA1},
{8'hAF, 8'hB7, 8'h88},
{8'hBF, 8'hC5, 8'hA3},
{8'hE6, 8'hE9, 8'hD4},
{8'hDC, 8'hDF, 8'hCA},
{8'hD2, 8'hD5, 8'hBF},
{8'hDF, 8'hE1, 8'hD6},
{8'hE1, 8'hE4, 8'hCF},
{8'hDE, 8'hE2, 8'hC4},
{8'hD0, 8'hD2, 8'hB9},
{8'hC4, 8'hC3, 8'hB3},
{8'hEF, 8'hED, 8'hDF},
{8'hE5, 8'hE4, 8'hCD},
{8'hDF, 8'hDE, 8'hC0},
{8'hC6, 8'hC7, 8'hB6},
{8'h97, 8'h99, 8'h80},
{8'hB0, 8'hB6, 8'h8E},
{8'hD7, 8'hDF, 8'hAE},
{8'hDC, 8'hE4, 8'hB6},
{8'hE0, 8'hE7, 8'hC6},
{8'hF3, 8'hF7, 8'hE9},
{8'hF8, 8'hFA, 8'hF7},
{8'hFC, 8'hF9, 8'hF5},
{8'hFF, 8'hFD, 8'hFA},
{8'hFF, 8'hFE, 8'hFA},
{8'hFC, 8'hFA, 8'hF4},
{8'hF3, 8'hF2, 8'hEA},
{8'hDD, 8'hDE, 8'hD3},
{8'hE8, 8'hEA, 8'hDE},
{8'hE6, 8'hEA, 8'hD9},
{8'hE0, 8'hF2, 8'hB8},
{8'hE2, 8'hF4, 8'hB7},
{8'hE1, 8'hF3, 8'hB8},
{8'hE1, 8'hF0, 8'hBD},
{8'hE9, 8'hF5, 8'hCE},
{8'hC8, 8'hD1, 8'hB9},
{8'h7B, 8'h80, 8'h76},
{8'h7C, 8'h7E, 8'h7D},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'h7E, 8'h79, 8'h8C},
{8'h80, 8'h7E, 8'h82},
{8'h9E, 8'h9F, 8'h8E},
{8'hBA, 8'hBD, 8'h9D},
{8'hC3, 8'hC7, 8'hA5},
{8'hA3, 8'hA4, 8'h8F},
{8'hA0, 8'h9F, 8'h9D},
{8'hDE, 8'hDC, 8'hE5},
{8'hF5, 8'hF6, 8'hF6},
{8'hFF, 8'hFF, 8'hFD},
{8'hFE, 8'hFF, 8'hFA},
{8'hF7, 8'hF7, 8'hEF},
{8'hF5, 8'hF4, 8'hEB},
{8'hF9, 8'hF5, 8'hEC},
{8'hFC, 8'hF8, 8'hEF},
{8'hFD, 8'hF9, 8'hEF},
{8'hF6, 8'hF5, 8'hDA},
{8'hEB, 8'hE9, 8'hCB},
{8'hE8, 8'hE5, 8'hC8},
{8'hEA, 8'hE7, 8'hCB},
{8'hE9, 8'hE7, 8'hD2},
{8'hEC, 8'hEA, 8'hE1},
{8'hF3, 8'hF0, 8'hF1},
{8'hF6, 8'hF3, 8'hF9},
{8'hF7, 8'hF4, 8'hF7},
{8'hF8, 8'hF5, 8'hF6},
{8'hF0, 8'hED, 8'hE2},
{8'hF3, 8'hF1, 8'hCE},
{8'hE7, 8'hE5, 8'hA9},
{8'hE5, 8'hE2, 8'h9B},
{8'hEB, 8'hE6, 8'hA3},
{8'hFB, 8'hF4, 8'hC0},
{8'hEE, 8'hED, 8'hE0},
{8'hF5, 8'hF5, 8'hEE},
{8'hFC, 8'hFB, 8'hF6},
{8'hF7, 8'hF6, 8'hF1},
{8'hF4, 8'hF4, 8'hED},
{8'hD9, 8'hD9, 8'hCE},
{8'hC6, 8'hC7, 8'hB7},
{8'hD3, 8'hD4, 8'hC1},
{8'hEA, 8'hE7, 8'hDF},
{8'hF0, 8'hF1, 8'hF1},
{8'hF7, 8'hFA, 8'hFF},
{8'hD7, 8'hD5, 8'hDE},
{8'h15, 8'h0F, 8'h19},
{8'h02, 8'h00, 8'h12},
{8'h00, 8'h00, 8'h23},
{8'h0F, 8'h20, 8'h52},
{8'h1C, 8'h51, 8'hA6},
{8'h0F, 8'h53, 8'hBB},
{8'h21, 8'h51, 8'hAE},
{8'h19, 8'h54, 8'hBB},
{8'h28, 8'h59, 8'hB3},
{8'h3E, 8'h53, 8'h8B},
{8'h10, 8'h29, 8'h59},
{8'h8B, 8'h91, 8'hA4},
{8'hF1, 8'hDB, 8'hE7},
{8'hDE, 8'hCC, 8'hD7},
{8'hED, 8'hE4, 8'hEB},
{8'hFF, 8'hFF, 8'hFF},
{8'hFE, 8'hFF, 8'hFF},
{8'hFC, 8'hFF, 8'hFF},
{8'hFE, 8'hFF, 8'hFF},
{8'hFE, 8'hFF, 8'hFD},
{8'hF9, 8'hFA, 8'hFA},
{8'hFF, 8'hFF, 8'hFF},
{8'hC5, 8'hC4, 8'hC9},
{8'h4D, 8'h48, 8'h61},
{8'h52, 8'h50, 8'h55},
{8'h81, 8'h7D, 8'h8A},
{8'hFC, 8'hFD, 8'hF6},
{8'hFB, 8'hFC, 8'hF3},
{8'hF7, 8'hF7, 8'hF4},
{8'hD3, 8'hD5, 8'hC7},
{8'hE5, 8'hE9, 8'hD1},
{8'hE0, 8'hE2, 8'hCF},
{8'hF1, 8'hF3, 8'hEA},
{8'hF0, 8'hF0, 8'hEC},
{8'hDB, 8'hDD, 8'hD3},
{8'hBA, 8'hBD, 8'hAA},
{8'hD0, 8'hD7, 8'hBC},
{8'hDF, 8'hE7, 8'hC4},
{8'hE6, 8'hEE, 8'hC5},
{8'hC3, 8'hC9, 8'hA9},
{8'hA3, 8'hA5, 8'h96},
{8'hD9, 8'hD9, 8'hD2},
{8'hEF, 8'hED, 8'hE2},
{8'hEB, 8'hEB, 8'hD7},
{8'hD4, 8'hDB, 8'hBD},
{8'hA3, 8'hAB, 8'h8A},
{8'hC1, 8'hC8, 8'hA4},
{8'hD3, 8'hDA, 8'hB3},
{8'hDC, 8'hE2, 8'hBD},
{8'hE8, 8'hEB, 8'hCD},
{8'hE7, 8'hE8, 8'hD1},
{8'hE2, 8'hE2, 8'hD1},
{8'hE0, 8'hDD, 8'hCE},
{8'hEA, 8'hE6, 8'hDD},
{8'hF1, 8'hEE, 8'hEB},
{8'hF0, 8'hEF, 8'hEF},
{8'hF0, 8'hEF, 8'hEE},
{8'hE7, 8'hE8, 8'hE0},
{8'hE2, 8'hE4, 8'hD3},
{8'hEA, 8'hEF, 8'hD5},
{8'hE2, 8'hF4, 8'hB9},
{8'hE1, 8'hF3, 8'hB7},
{8'hE1, 8'hF1, 8'hBA},
{8'hE1, 8'hEE, 8'hC1},
{8'hE8, 8'hF2, 8'hD1},
{8'hAB, 8'hB2, 8'hA0},
{8'h79, 8'h7C, 8'h77},
{8'h7D, 8'h7D, 8'h81},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'h7F, 8'h79, 8'h94},
{8'h82, 8'h7F, 8'h88},
{8'h78, 8'h79, 8'h66},
{8'hBC, 8'hC1, 8'h98},
{8'hF4, 8'hFA, 8'hCB},
{8'hEF, 8'hF3, 8'hD0},
{8'hE8, 8'hE8, 8'hDA},
{8'hF4, 8'hF3, 8'hF1},
{8'hF3, 8'hF5, 8'hEA},
{8'hF6, 8'hF7, 8'hED},
{8'hF4, 8'hF5, 8'hEC},
{8'hEE, 8'hEE, 8'hE6},
{8'hF3, 8'hF2, 8'hEA},
{8'hF5, 8'hF2, 8'hE8},
{8'hF5, 8'hF2, 8'hE5},
{8'hF6, 8'hF2, 8'hE2},
{8'hF0, 8'hEE, 8'hC7},
{8'hE8, 8'hE7, 8'hC2},
{8'hDE, 8'hDE, 8'hC0},
{8'hEC, 8'hEE, 8'hD8},
{8'hE7, 8'hE9, 8'hDC},
{8'hEF, 8'hF0, 8'hED},
{8'hEF, 8'hEF, 8'hF3},
{8'hF7, 8'hF5, 8'hFD},
{8'hF9, 8'hF3, 8'hF6},
{8'hFE, 8'hF8, 8'hF8},
{8'hF7, 8'hEF, 8'hE5},
{8'hF5, 8'hF0, 8'hCC},
{8'hE8, 8'hE6, 8'hA5},
{8'hD4, 8'hD2, 8'h81},
{8'hE0, 8'hDB, 8'h8B},
{8'hFA, 8'hF5, 8'hB2},
{8'hF1, 8'hF0, 8'hE4},
{8'hF7, 8'hF6, 8'hF2},
{8'hFB, 8'hFA, 8'hF8},
{8'hFA, 8'hF9, 8'hF8},
{8'hF5, 8'hF4, 8'hF3},
{8'hFE, 8'hFD, 8'hF8},
{8'hF5, 8'hF6, 8'hEB},
{8'hD9, 8'hD9, 8'hCC},
{8'hEC, 8'hE8, 8'hE6},
{8'hF6, 8'hF7, 8'hF7},
{8'hF2, 8'hF5, 8'hF5},
{8'hDC, 8'hDB, 8'hDA},
{8'h1A, 8'h16, 8'h1A},
{8'h01, 8'h02, 8'h18},
{8'h01, 8'h08, 8'h3B},
{8'h1E, 8'h3E, 8'h87},
{8'h0E, 8'h56, 8'hBC},
{8'h03, 8'h52, 8'hC3},
{8'h1D, 8'h4E, 8'hAA},
{8'h20, 8'h52, 8'hAF},
{8'h32, 8'h56, 8'hA5},
{8'h85, 8'h91, 8'hC2},
{8'h28, 8'h42, 8'h74},
{8'h7F, 8'h86, 8'hA2},
{8'hE9, 8'hCE, 8'hD7},
{8'hE4, 8'hCD, 8'hD3},
{8'hF0, 8'hE4, 8'hE8},
{8'hFF, 8'hFD, 8'hFE},
{8'hFF, 8'hFF, 8'hFF},
{8'hFD, 8'hFF, 8'hFF},
{8'hFC, 8'hFF, 8'hFF},
{8'hFD, 8'hFF, 8'hFD},
{8'hFE, 8'hFD, 8'hF7},
{8'hF4, 8'hF2, 8'hF5},
{8'hEF, 8'hF0, 8'hEF},
{8'h5E, 8'h5C, 8'h7A},
{8'h25, 8'h27, 8'h29},
{8'h11, 8'h10, 8'h23},
{8'hBE, 8'hC1, 8'hB9},
{8'hFC, 8'hFD, 8'hF5},
{8'hF7, 8'hF7, 8'hF2},
{8'hF2, 8'hF4, 8'hE8},
{8'hF8, 8'hF9, 8'hEE},
{8'hFE, 8'hFE, 8'hFD},
{8'hFC, 8'hF9, 8'hFF},
{8'hFF, 8'hFE, 8'hFF},
{8'hF6, 8'hF7, 8'hF0},
{8'hC7, 8'hCB, 8'hB3},
{8'hD2, 8'hDF, 8'hB1},
{8'hEA, 8'hF8, 8'hC2},
{8'hE3, 8'hF0, 8'hBB},
{8'hBC, 8'hC4, 8'h9D},
{8'h89, 8'h8D, 8'h7D},
{8'hC2, 8'hC2, 8'hC1},
{8'hF5, 8'hF4, 8'hF3},
{8'hF7, 8'hF8, 8'hEF},
{8'hBC, 8'hCA, 8'hA7},
{8'h97, 8'hA4, 8'h84},
{8'hD8, 8'hE1, 8'hC8},
{8'hDF, 8'hE2, 8'hD0},
{8'hF5, 8'hF6, 8'hE5},
{8'hFD, 8'hFD, 8'hEA},
{8'hF7, 8'hF5, 8'hE0},
{8'hDF, 8'hDB, 8'hC2},
{8'hE1, 8'hDF, 8'hC7},
{8'hEE, 8'hEA, 8'hDC},
{8'hF7, 8'hF3, 8'hF2},
{8'hF9, 8'hF6, 8'hF9},
{8'hFB, 8'hF9, 8'hFD},
{8'hEE, 8'hEF, 8'hE7},
{8'hDD, 8'hE0, 8'hCA},
{8'hE1, 8'hE8, 8'hC4},
{8'hE1, 8'hF2, 8'hB9},
{8'hE2, 8'hF3, 8'hBA},
{8'hE5, 8'hF3, 8'hC3},
{8'hE6, 8'hF1, 8'hCB},
{8'hB8, 8'hC0, 8'hA8},
{8'h7C, 8'h80, 8'h76},
{8'h82, 8'h83, 8'h85},
{8'h7A, 8'h79, 8'h83},
{8'h7F, 8'h7D, 8'h81},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'h7D, 8'h7B, 8'h84},
{8'h7D, 8'h7B, 8'h7D},
{8'h78, 8'h78, 8'h6E},
{8'h8D, 8'h8F, 8'h78},
{8'hE9, 8'hEC, 8'hCC},
{8'hF0, 8'hF5, 8'hD1},
{8'hEB, 8'hEF, 8'hCC},
{8'hEE, 8'hF2, 8'hD1},
{8'hE7, 8'hEC, 8'hD3},
{8'hEB, 8'hEE, 8'hDB},
{8'hEE, 8'hEF, 8'hE4},
{8'hF5, 8'hF4, 8'hF0},
{8'hFD, 8'hFB, 8'hF6},
{8'hFB, 8'hF9, 8'hEE},
{8'hF8, 8'hF5, 8'hE3},
{8'hF5, 8'hF3, 8'hDB},
{8'hF6, 8'hF0, 8'hCA},
{8'hEC, 8'hE8, 8'hC6},
{8'hE4, 8'hE2, 8'hCB},
{8'hF0, 8'hF2, 8'hE4},
{8'hE5, 8'hE9, 8'hE0},
{8'hB8, 8'hBC, 8'hB3},
{8'hA7, 8'hA9, 8'h9E},
{8'hBE, 8'hC0, 8'hB2},
{8'hF6, 8'hEF, 8'hE9},
{8'hFA, 8'hF1, 8'hEE},
{8'hF9, 8'hF0, 8'hE8},
{8'hF6, 8'hEE, 8'hD5},
{8'hF3, 8'hED, 8'hBE},
{8'hDE, 8'hD9, 8'h9F},
{8'hE6, 8'hDF, 8'hA8},
{8'hF9, 8'hF2, 8'hC6},
{8'hF1, 8'hF0, 8'hE5},
{8'hF6, 8'hF5, 8'hEF},
{8'hFB, 8'hFB, 8'hF8},
{8'hF3, 8'hF2, 8'hF1},
{8'hFE, 8'hFD, 8'hFC},
{8'hF9, 8'hF8, 8'hF5},
{8'hFB, 8'hFB, 8'hF4},
{8'hEF, 8'hEE, 8'hE5},
{8'hF4, 8'hF0, 8'hEE},
{8'hF1, 8'hF1, 8'hEE},
{8'hF7, 8'hFA, 8'hF5},
{8'hC0, 8'hC0, 8'hBA},
{8'h07, 8'h06, 8'h08},
{8'h00, 8'h01, 8'h1E},
{8'h0D, 8'h21, 8'h63},
{8'h22, 8'h4E, 8'hAA},
{8'h0B, 8'h58, 8'hC5},
{8'h06, 8'h5A, 8'hCD},
{8'h1D, 8'h4E, 8'hA9},
{8'h1D, 8'h51, 8'hAD},
{8'h28, 8'h53, 8'hA6},
{8'h5A, 8'h76, 8'hB5},
{8'h1C, 8'h4E, 8'h98},
{8'h4B, 8'h6C, 8'hA6},
{8'hDC, 8'hC3, 8'hCD},
{8'hE5, 8'hCD, 8'hD2},
{8'hFB, 8'hF0, 8'hF4},
{8'hFC, 8'hF9, 8'hFA},
{8'hFF, 8'hFE, 8'hFF},
{8'hFD, 8'hFF, 8'hFF},
{8'hFC, 8'hFF, 8'hFF},
{8'hFD, 8'hFF, 8'hFE},
{8'hFE, 8'hFD, 8'hF7},
{8'hEC, 8'hE9, 8'hEC},
{8'hEA, 8'hEB, 8'hF3},
{8'h9F, 8'hA1, 8'hB4},
{8'h06, 8'h08, 8'h1B},
{8'h00, 8'h00, 8'h0E},
{8'h37, 8'h37, 8'h3C},
{8'hE0, 8'hE1, 8'hDE},
{8'hF2, 8'hF4, 8'hE3},
{8'hF9, 8'hFA, 8'hE7},
{8'hF9, 8'hF9, 8'hEB},
{8'hFA, 8'hF9, 8'hF7},
{8'hFA, 8'hF7, 8'hFD},
{8'hFE, 8'hFC, 8'hFE},
{8'hED, 8'hEE, 8'hDF},
{8'hC2, 8'hC6, 8'hA2},
{8'hD2, 8'hE1, 8'hA6},
{8'hE5, 8'hF4, 8'hB4},
{8'hE1, 8'hF0, 8'hB1},
{8'hCB, 8'hD6, 8'hAB},
{8'h8E, 8'h92, 8'h82},
{8'hCC, 8'hCD, 8'hCE},
{8'hF6, 8'hF5, 8'hFB},
{8'hF7, 8'hF8, 8'hF7},
{8'hCA, 8'hD8, 8'hBE},
{8'hC2, 8'hCF, 8'hBC},
{8'hE4, 8'hEB, 8'hE6},
{8'hFA, 8'hFC, 8'hFE},
{8'hFB, 8'hF8, 8'hFB},
{8'hFA, 8'hF3, 8'hF2},
{8'hFF, 8'hFB, 8'hEF},
{8'hEA, 8'hE4, 8'hCF},
{8'hE1, 8'hDF, 8'hC0},
{8'hE5, 8'hE3, 8'hCE},
{8'hF2, 8'hEE, 8'hE8},
{8'hF6, 8'hF3, 8'hF6},
{8'hF6, 8'hF4, 8'hF6},
{8'hF1, 8'hF3, 8'hE7},
{8'hE6, 8'hEB, 8'hCE},
{8'hE4, 8'hEB, 8'hC2},
{8'hE5, 8'hF2, 8'hC0},
{8'hDC, 8'hE9, 8'hBA},
{8'hBF, 8'hCA, 8'hA3},
{8'hC6, 8'hCE, 8'hB3},
{8'h7E, 8'h82, 8'h73},
{8'h7E, 8'h7F, 8'h7D},
{8'h7D, 8'h7B, 8'h82},
{8'h82, 8'h7F, 8'h8B},
{8'h80, 8'h7E, 8'h82},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'h7D, 8'h7D, 8'h70},
{8'h7F, 8'h7F, 8'h77},
{8'h80, 8'h7F, 8'h7E},
{8'h7C, 8'h7B, 8'h7B},
{8'hBC, 8'hBC, 8'hB2},
{8'hF5, 8'hF8, 8'hDC},
{8'hEA, 8'hF1, 8'hBE},
{8'hE7, 8'hF0, 8'hB2},
{8'hCD, 8'hD5, 8'hAD},
{8'hEA, 8'hEE, 8'hD2},
{8'hF4, 8'hF6, 8'hE8},
{8'hFA, 8'hF9, 8'hF5},
{8'hFE, 8'hFC, 8'hF9},
{8'hFC, 8'hF9, 8'hEE},
{8'hF7, 8'hF5, 8'hDF},
{8'hF3, 8'hF2, 8'hD3},
{8'hFC, 8'hF0, 8'hC2},
{8'hF5, 8'hEC, 8'hC5},
{8'hE6, 8'hE3, 8'hCB},
{8'hE1, 8'hE3, 8'hD5},
{8'h88, 8'h8E, 8'h81},
{8'h7C, 8'h83, 8'h6E},
{8'h96, 8'h9C, 8'h7B},
{8'hB3, 8'hB7, 8'h8F},
{8'hF6, 8'hF1, 8'hDD},
{8'hF9, 8'hF1, 8'hE8},
{8'hF7, 8'hEE, 8'hEA},
{8'hFB, 8'hF3, 8'hE9},
{8'hFB, 8'hF5, 8'hDE},
{8'hEE, 8'hE8, 8'hCE},
{8'hF7, 8'hF0, 8'hDF},
{8'hF8, 8'hF0, 8'hE8},
{8'hF1, 8'hF2, 8'hE2},
{8'hED, 8'hEE, 8'hDF},
{8'hFA, 8'hFA, 8'hF1},
{8'hF6, 8'hF6, 8'hF0},
{8'hF8, 8'hF7, 8'hF2},
{8'hFC, 8'hFC, 8'hF6},
{8'hFE, 8'hFE, 8'hF4},
{8'hD2, 8'hD2, 8'hC6},
{8'hEB, 8'hE7, 8'hDD},
{8'hF7, 8'hF7, 8'hEE},
{8'hF8, 8'hFB, 8'hF3},
{8'h97, 8'h97, 8'h92},
{8'h01, 8'h01, 8'h06},
{8'h00, 8'h01, 8'h28},
{8'h16, 8'h37, 8'h84},
{8'h1B, 8'h50, 8'hB7},
{8'h0F, 8'h54, 8'hBD},
{8'h07, 8'h56, 8'hC5},
{8'h1D, 8'h50, 8'hAA},
{8'h15, 8'h52, 8'hB3},
{8'h18, 8'h54, 8'hB2},
{8'h1B, 8'h4C, 8'hA0},
{8'h0A, 8'h58, 8'hBD},
{8'h1F, 8'h5E, 8'hB4},
{8'hCD, 8'hBC, 8'hCD},
{8'hEB, 8'hD8, 8'hE2},
{8'hFE, 8'hF7, 8'hFD},
{8'hFD, 8'hFB, 8'hFD},
{8'hFE, 8'hFF, 8'hFF},
{8'hFD, 8'hFF, 8'hFF},
{8'hFE, 8'hFF, 8'hFF},
{8'hFE, 8'hFE, 8'hFF},
{8'hFE, 8'hF9, 8'hF4},
{8'hF7, 8'hF5, 8'hF2},
{8'hD4, 8'hD3, 8'hF0},
{8'hC7, 8'hCE, 8'hDE},
{8'h1D, 8'h22, 8'h4E},
{8'h00, 8'h04, 8'h13},
{8'h00, 8'h00, 8'h13},
{8'h57, 8'h58, 8'h5D},
{8'hF4, 8'hF5, 8'hDC},
{8'hF4, 8'hF4, 8'hD8},
{8'hF9, 8'hFA, 8'hE0},
{8'hF9, 8'hF8, 8'hE8},
{8'hFB, 8'hF9, 8'hF4},
{8'hF5, 8'hF3, 8'hEC},
{8'hE7, 8'hE7, 8'hCF},
{8'hD1, 8'hD4, 8'hAA},
{8'hD3, 8'hE0, 8'hA1},
{8'hE8, 8'hF6, 8'hB2},
{8'hD7, 8'hE3, 8'hA2},
{8'hC6, 8'hCE, 8'hA0},
{8'hB7, 8'hB9, 8'hA7},
{8'hEF, 8'hED, 8'hED},
{8'hFA, 8'hF7, 8'hFC},
{8'hF4, 8'hF2, 8'hF2},
{8'hEC, 8'hF5, 8'hE9},
{8'hB1, 8'hBA, 8'hB4},
{8'hF1, 8'hF6, 8'hF7},
{8'hF8, 8'hF7, 8'hFF},
{8'hFD, 8'hF9, 8'hFF},
{8'hFB, 8'hF5, 8'hFB},
{8'hFE, 8'hFA, 8'hF6},
{8'hE5, 8'hDF, 8'hD1},
{8'hD7, 8'hD6, 8'hB5},
{8'hDC, 8'hDB, 8'hBF},
{8'hE4, 8'hE3, 8'hD1},
{8'hF2, 8'hF1, 8'hE6},
{8'hEA, 8'hEB, 8'hDE},
{8'hF3, 8'hF6, 8'hE0},
{8'hF2, 8'hF7, 8'hD4},
{8'hE8, 8'hF0, 8'hC5},
{8'hDC, 8'hE7, 8'hBF},
{8'h9F, 8'hA9, 8'h87},
{8'h83, 8'h8A, 8'h70},
{8'h84, 8'h88, 8'h79},
{8'h7D, 8'h7E, 8'h79},
{8'h7E, 8'h7E, 8'h80},
{8'h7F, 8'h7C, 8'h84},
{8'h7F, 8'h7C, 8'h85},
{8'h7F, 8'h7D, 8'h81},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'h7E, 8'h7E, 8'h71},
{8'h7D, 8'h7C, 8'h76},
{8'h7E, 8'h7D, 8'h7D},
{8'h7E, 8'h7C, 8'h7D},
{8'h7C, 8'h7C, 8'h74},
{8'hB8, 8'hBB, 8'hA0},
{8'hE9, 8'hEF, 8'hBE},
{8'hE8, 8'hF0, 8'hB3},
{8'hC9, 8'hD2, 8'hA0},
{8'hEB, 8'hF1, 8'hCD},
{8'hF2, 8'hF5, 8'hE3},
{8'hF4, 8'hF3, 8'hEF},
{8'hFD, 8'hFA, 8'hF8},
{8'hF9, 8'hF6, 8'hEB},
{8'hF4, 8'hF2, 8'hD9},
{8'hF2, 8'hF1, 8'hCA},
{8'hF8, 8'hEB, 8'h9E},
{8'hF2, 8'hE5, 8'hA4},
{8'hF5, 8'hF0, 8'hC7},
{8'hE5, 8'hE6, 8'hD1},
{8'h9D, 8'hA1, 8'h92},
{8'h86, 8'h89, 8'h74},
{8'hAA, 8'hAC, 8'h88},
{8'hA2, 8'hA2, 8'h75},
{8'hF2, 8'hEF, 8'hDB},
{8'hFB, 8'hF6, 8'hF0},
{8'hF9, 8'hF4, 8'hF5},
{8'hFC, 8'hF7, 8'hF6},
{8'hF5, 8'hF1, 8'hE8},
{8'hF4, 8'hF2, 8'hE6},
{8'hFC, 8'hF9, 8'hF6},
{8'hDA, 8'hD5, 8'hDB},
{8'hBB, 8'hBE, 8'hA4},
{8'hD1, 8'hD3, 8'hB9},
{8'hF3, 8'hF4, 8'hE1},
{8'hF0, 8'hF1, 8'hE2},
{8'hEC, 8'hED, 8'hDF},
{8'hF1, 8'hF2, 8'hE4},
{8'hF6, 8'hF7, 8'hE6},
{8'hEE, 8'hEF, 8'hDB},
{8'hF0, 8'hED, 8'hD5},
{8'hF5, 8'hF6, 8'hE5},
{8'hE6, 8'hE8, 8'hE1},
{8'h34, 8'h32, 8'h37},
{8'h00, 8'h00, 8'h13},
{8'h02, 8'h05, 8'h36},
{8'h1B, 8'h46, 8'h99},
{8'h11, 8'h51, 8'hBA},
{8'h15, 8'h52, 8'hB6},
{8'h0B, 8'h55, 8'hC0},
{8'h1C, 8'h50, 8'hAB},
{8'h11, 8'h55, 8'hBA},
{8'h10, 8'h55, 8'hBB},
{8'h17, 8'h50, 8'hAB},
{8'h07, 8'h56, 8'hC3},
{8'h0B, 8'h4A, 8'hA7},
{8'h84, 8'h7C, 8'h95},
{8'hE1, 8'hD8, 8'hE8},
{8'hFF, 8'hFF, 8'hFF},
{8'hFA, 8'hFD, 8'hFF},
{8'hFB, 8'hFF, 8'hFF},
{8'hFD, 8'hFF, 8'hFF},
{8'hFF, 8'hFF, 8'hFD},
{8'hFF, 8'hFE, 8'hFD},
{8'hFF, 8'hFA, 8'hF7},
{8'hFB, 8'hF5, 8'hF4},
{8'hD4, 8'hD2, 8'hF4},
{8'h84, 8'h8B, 8'hA7},
{8'h13, 8'h18, 8'h4D},
{8'h05, 8'h0B, 8'h26},
{8'h04, 8'h07, 8'h25},
{8'h00, 8'h00, 8'h0E},
{8'h81, 8'h7F, 8'h70},
{8'hF0, 8'hEF, 8'hD5},
{8'hFD, 8'hFE, 8'hE0},
{8'hFA, 8'hF9, 8'hDE},
{8'hF8, 8'hF6, 8'hE5},
{8'hED, 8'hEB, 8'hDC},
{8'hDE, 8'hDC, 8'hC6},
{8'hCB, 8'hCC, 8'hA9},
{8'hD9, 8'hE1, 8'hA7},
{8'hE2, 8'hEB, 8'hAC},
{8'hD4, 8'hDB, 8'h9E},
{8'hCC, 8'hCF, 8'hA2},
{8'hBD, 8'hBB, 8'hA6},
{8'hF7, 8'hF1, 8'hED},
{8'hFB, 8'hF4, 8'hF2},
{8'hF9, 8'hF3, 8'hEC},
{8'hEF, 8'hF2, 8'hEC},
{8'hC7, 8'hCB, 8'hC6},
{8'hFE, 8'hFF, 8'hFD},
{8'hFC, 8'hFC, 8'hFB},
{8'hF9, 8'hF9, 8'hF9},
{8'hF7, 8'hF5, 8'hF0},
{8'hF5, 8'hF4, 8'hEA},
{8'hD2, 8'hD1, 8'hC1},
{8'hCD, 8'hCC, 8'hAE},
{8'hDC, 8'hDC, 8'hBD},
{8'hE1, 8'hE2, 8'hC1},
{8'hE6, 8'hE9, 8'hC8},
{8'hD7, 8'hDB, 8'hB7},
{8'hDB, 8'hE2, 8'hBC},
{8'hDD, 8'hE3, 8'hBB},
{8'hD1, 8'hD9, 8'hB1},
{8'hA4, 8'hAD, 8'h92},
{8'h89, 8'h8F, 8'h7B},
{8'h7E, 8'h81, 8'h76},
{8'h81, 8'h81, 8'h7F},
{8'h7F, 8'h7E, 8'h80},
{8'h7F, 8'h7D, 8'h82},
{8'h7F, 8'h7D, 8'h81},
{8'h81, 8'h7C, 8'h80},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'h84, 8'h81, 8'h89},
{8'h88, 8'h86, 8'h88},
{8'h90, 8'h90, 8'h87},
{8'h96, 8'h97, 8'h83},
{8'h9B, 8'h9E, 8'h82},
{8'h92, 8'h96, 8'h75},
{8'h94, 8'h98, 8'h75},
{8'hD8, 8'hDD, 8'hB7},
{8'hC1, 8'hCB, 8'h94},
{8'hE6, 8'hEE, 8'hC4},
{8'hF0, 8'hF3, 8'hE0},
{8'hF6, 8'hF6, 8'hF4},
{8'hFE, 8'hFC, 8'hFD},
{8'hFD, 8'hFA, 8'hEF},
{8'hF7, 8'hF7, 8'hDB},
{8'hF6, 8'hF5, 8'hC5},
{8'hEC, 8'hDC, 8'h61},
{8'hE0, 8'hD2, 8'h67},
{8'hF0, 8'hEA, 8'hA6},
{8'hFD, 8'hFD, 8'hDC},
{8'hF5, 8'hF8, 8'hEA},
{8'hC4, 8'hC4, 8'hB7},
{8'hB9, 8'hB5, 8'h9F},
{8'hC6, 8'hC1, 8'hA4},
{8'hF8, 8'hF6, 8'hEC},
{8'hF3, 8'hEF, 8'hF2},
{8'hFB, 8'hF8, 8'hFF},
{8'hF7, 8'hF5, 8'hF9},
{8'hF9, 8'hFA, 8'hF0},
{8'hF7, 8'hFA, 8'hE7},
{8'hFA, 8'hFE, 8'hEF},
{8'hCF, 8'hD1, 8'hC7},
{8'hA5, 8'hAA, 8'h84},
{8'hC3, 8'hC7, 8'hA2},
{8'hC3, 8'hC7, 8'hA7},
{8'hE0, 8'hE3, 8'hC8},
{8'hF0, 8'hF2, 8'hDA},
{8'hEB, 8'hED, 8'hD5},
{8'hF1, 8'hF4, 8'hDA},
{8'hED, 8'hEF, 8'hD4},
{8'hED, 8'hED, 8'hC8},
{8'hEC, 8'hED, 8'hD3},
{8'h90, 8'h91, 8'h8B},
{8'h02, 8'h01, 8'h0D},
{8'h02, 8'h00, 8'h23},
{8'h05, 8'h11, 8'h4B},
{8'h19, 8'h4B, 8'hA1},
{8'h0F, 8'h56, 8'hBE},
{8'h18, 8'h51, 8'hB4},
{8'h0C, 8'h54, 8'hBF},
{8'h1A, 8'h51, 8'hAC},
{8'h0D, 8'h56, 8'hBD},
{8'h10, 8'h56, 8'hBB},
{8'h16, 8'h45, 8'h99},
{8'h10, 8'h4E, 8'hAE},
{8'h1F, 8'h45, 8'h96},
{8'h07, 8'h07, 8'h25},
{8'h3C, 8'h3C, 8'h54},
{8'hB5, 8'hB9, 8'hC6},
{8'hF3, 8'hF9, 8'hFB},
{8'hFF, 8'hFF, 8'hFF},
{8'hFF, 8'hFF, 8'hFF},
{8'hFF, 8'hFF, 8'hFC},
{8'hFF, 8'hFE, 8'hF9},
{8'hFF, 8'hF9, 8'hF8},
{8'hFF, 8'hF6, 8'hFE},
{8'hC3, 8'hC2, 8'hDA},
{8'h3C, 8'h42, 8'h74},
{8'h05, 8'h0E, 8'h3D},
{8'h0A, 8'h0F, 8'h3F},
{8'h04, 8'h05, 8'h24},
{8'h04, 8'h04, 8'h1D},
{8'h0D, 8'h07, 8'h0A},
{8'hA7, 8'hA4, 8'h94},
{8'hFF, 8'hFF, 8'hE4},
{8'hF2, 8'hF2, 8'hD3},
{8'hF1, 8'hEE, 8'hD9},
{8'hF8, 8'hF5, 8'hE9},
{8'hF8, 8'hF5, 8'hEA},
{8'hE4, 8'hE1, 8'hD0},
{8'hDE, 8'hE1, 8'hB1},
{8'hDD, 8'hE0, 8'hA7},
{8'hD2, 8'hD4, 8'h9A},
{8'hD1, 8'hD0, 8'hA3},
{8'hE2, 8'hDC, 8'hC4},
{8'hFB, 8'hF3, 8'hEA},
{8'hFB, 8'hF1, 8'hE8},
{8'hF8, 8'hEF, 8'hDF},
{8'hEC, 8'hEC, 8'hE1},
{8'hE3, 8'hE5, 8'hD7},
{8'hF7, 8'hFA, 8'hE7},
{8'hEB, 8'hEF, 8'hD6},
{8'hEC, 8'hF0, 8'hD5},
{8'hF0, 8'hF4, 8'hD9},
{8'hE1, 8'hE6, 8'hCB},
{8'hB6, 8'hBC, 8'hA2},
{8'hB4, 8'hB3, 8'h9A},
{8'hCF, 8'hCE, 8'hAD},
{8'hD5, 8'hD8, 8'hAA},
{8'hD8, 8'hDD, 8'hA6},
{8'hD8, 8'hE1, 8'hA7},
{8'hCA, 8'hD3, 8'h9D},
{8'hD1, 8'hD8, 8'hAB},
{8'hAB, 8'hB2, 8'h8E},
{8'h7A, 8'h7E, 8'h70},
{8'h7D, 8'h80, 8'h77},
{8'h7F, 8'h81, 8'h7F},
{8'h7D, 8'h7D, 8'h82},
{8'h7E, 8'h7C, 8'h83},
{8'h7F, 8'h7D, 8'h81},
{8'h81, 8'h7D, 8'h7D},
{8'h81, 8'h7D, 8'h7A},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'h80, 8'h7D, 8'h89},
{8'h81, 8'h7F, 8'h84},
{8'h81, 8'h81, 8'h79},
{8'h82, 8'h83, 8'h6F},
{8'hD2, 8'hD5, 8'hBA},
{8'hD4, 8'hD7, 8'hBA},
{8'hC1, 8'hC4, 8'hA9},
{8'hD8, 8'hDB, 8'hBF},
{8'hB1, 8'hB6, 8'h84},
{8'hEE, 8'hF2, 8'hC9},
{8'hFC, 8'hFC, 8'hE7},
{8'hFC, 8'hFA, 8'hF1},
{8'hFE, 8'hFD, 8'hF7},
{8'hFE, 8'hFD, 8'hEF},
{8'hFA, 8'hFB, 8'hDF},
{8'hF6, 8'hF8, 8'hCE},
{8'hE6, 8'hDD, 8'h79},
{8'hD9, 8'hD1, 8'h79},
{8'hEA, 8'hE6, 8'hAB},
{8'hFA, 8'hF8, 8'hD8},
{8'hF8, 8'hF6, 8'hE7},
{8'hDB, 8'hD8, 8'hCC},
{8'hC2, 8'hBC, 8'hAC},
{8'hF4, 8'hF0, 8'hDB},
{8'hF1, 8'hF0, 8'hE5},
{8'hF3, 8'hF2, 8'hEE},
{8'hD5, 8'hD4, 8'hD4},
{8'hF0, 8'hEF, 8'hEC},
{8'hF9, 8'hFB, 8'hF1},
{8'hF6, 8'hF8, 8'hEA},
{8'hF8, 8'hFA, 8'hEE},
{8'hDF, 8'hE2, 8'hD6},
{8'hAA, 8'hAD, 8'h88},
{8'hC4, 8'hC6, 8'hA6},
{8'hDC, 8'hDC, 8'hC6},
{8'hEB, 8'hEB, 8'hDC},
{8'hFF, 8'hFC, 8'hF0},
{8'hFC, 8'hFC, 8'hE8},
{8'hF4, 8'hF5, 8'hD8},
{8'hE2, 8'hE5, 8'hBE},
{8'hDD, 8'hE2, 8'hA5},
{8'hD7, 8'hD7, 8'hBE},
{8'h2F, 8'h2B, 8'h35},
{8'h00, 8'h00, 8'h0F},
{8'h00, 8'h01, 8'h1F},
{8'h0D, 8'h1F, 8'h59},
{8'h18, 8'h4C, 8'hA5},
{8'h0F, 8'h55, 8'hBC},
{8'h10, 8'h55, 8'hAE},
{8'h0F, 8'h57, 8'hC5},
{8'h16, 8'h4E, 8'hB8},
{8'h19, 8'h55, 8'hB7},
{8'h0E, 8'h41, 8'h9E},
{8'h0D, 8'h30, 8'h8A},
{8'h1E, 8'h4E, 8'hA8},
{8'h1E, 8'h47, 8'h84},
{8'h08, 8'h08, 8'h2C},
{8'h00, 8'h00, 8'h18},
{8'h0E, 8'h10, 8'h3A},
{8'h62, 8'h73, 8'h9F},
{8'hA8, 8'hC4, 8'hD7},
{8'hE2, 8'hF9, 8'hFB},
{8'hFE, 8'hFF, 8'hFF},
{8'hFF, 8'hFF, 8'hF1},
{8'hFF, 8'hFC, 8'hF8},
{8'hEA, 8'hED, 8'hFC},
{8'h63, 8'h76, 8'hA2},
{8'h21, 8'h2F, 8'h72},
{8'h06, 8'h0A, 8'h2F},
{8'h09, 8'h13, 8'h41},
{8'h04, 8'h0C, 8'h27},
{8'h08, 8'h05, 8'h15},
{8'h02, 8'h00, 8'h13},
{8'h2C, 8'h27, 8'h28},
{8'hD9, 8'hD9, 8'hBB},
{8'hF0, 8'hF1, 8'hCA},
{8'hEC, 8'hEC, 8'hD1},
{8'hF8, 8'hF5, 8'hE9},
{8'hF8, 8'hF5, 8'hED},
{8'hF4, 8'hF1, 8'hE3},
{8'hDD, 8'hDF, 8'hB4},
{8'hD3, 8'hD4, 8'hA8},
{8'hD5, 8'hD3, 8'hAD},
{8'hF2, 8'hF0, 8'hD6},
{8'hF9, 8'hF2, 8'hE4},
{8'hFB, 8'hF4, 8'hEB},
{8'hFA, 8'hF1, 8'hE3},
{8'hF5, 8'hEC, 8'hD6},
{8'hF7, 8'hF1, 8'hD6},
{8'hF2, 8'hEF, 8'hD9},
{8'hF0, 8'hF0, 8'hDE},
{8'hF0, 8'hF4, 8'hDF},
{8'hF4, 8'hFA, 8'hE1},
{8'hE2, 8'hE9, 8'hCF},
{8'hE9, 8'hED, 8'hD9},
{8'hCE, 8'hD2, 8'hBF},
{8'hCA, 8'hCC, 8'hAE},
{8'hE4, 8'hE7, 8'hBF},
{8'hE6, 8'hEC, 8'hB8},
{8'hE8, 8'hF0, 8'hB7},
{8'hC6, 8'hCE, 8'h99},
{8'h9B, 8'hA2, 8'h7B},
{8'h9E, 8'hA1, 8'h8C},
{8'h82, 8'h84, 8'h7A},
{8'h7C, 8'h7D, 8'h77},
{8'h82, 8'h83, 8'h7F},
{8'h7E, 8'h7E, 8'h7F},
{8'h7E, 8'h7D, 8'h81},
{8'h7E, 8'h7C, 8'h81},
{8'h81, 8'h7E, 8'h82},
{8'h82, 8'h7F, 8'h80},
{8'h7E, 8'h7C, 8'h7B},
{8'h7F, 8'h7D, 8'h7F},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'h7F, 8'h7E, 8'h7F},
{8'h7D, 8'h7B, 8'h7E},
{8'h7E, 8'h7C, 8'h7E},
{8'h7B, 8'h79, 8'h78},
{8'hC1, 8'hC1, 8'hB8},
{8'hFD, 8'hFD, 8'hED},
{8'hE1, 8'hE3, 8'hC8},
{8'hC8, 8'hCB, 8'hAA},
{8'hC0, 8'hBC, 8'h9C},
{8'hF2, 8'hEE, 8'hD3},
{8'hF4, 8'hF0, 8'hDE},
{8'hF5, 8'hF1, 8'hE3},
{8'hFD, 8'hFA, 8'hEC},
{8'hF8, 8'hF8, 8'hE5},
{8'hF1, 8'hF5, 8'hDB},
{8'hED, 8'hF0, 8'hD0},
{8'hE6, 8'hE5, 8'hBE},
{8'hEA, 8'hE8, 8'hC5},
{8'hEE, 8'hEA, 8'hCE},
{8'hED, 8'hE9, 8'hD3},
{8'hEB, 8'hE6, 8'hD2},
{8'hD0, 8'hCB, 8'hB6},
{8'hD4, 8'hCF, 8'hB7},
{8'hF1, 8'hED, 8'hD2},
{8'hEE, 8'hEE, 8'hDA},
{8'hDD, 8'hDE, 8'hCB},
{8'hA0, 8'hA1, 8'h91},
{8'hD7, 8'hD7, 8'hCB},
{8'hFF, 8'hFF, 8'hF9},
{8'hF8, 8'hF7, 8'hF4},
{8'hF6, 8'hF4, 8'hF4},
{8'hEB, 8'hE9, 8'hE8},
{8'hC0, 8'hBF, 8'hA5},
{8'hEB, 8'hE8, 8'hD7},
{8'hFB, 8'hF7, 8'hF3},
{8'hFF, 8'hFD, 8'hFF},
{8'hFF, 8'hFC, 8'hFD},
{8'hFE, 8'hFA, 8'hEE},
{8'hF6, 8'hF5, 8'hD7},
{8'hE0, 8'hE3, 8'hB2},
{8'hDD, 8'hE7, 8'h97},
{8'h83, 8'h82, 8'h71},
{8'h05, 8'h00, 8'h1A},
{8'h07, 8'h03, 8'h1C},
{8'h00, 8'h03, 8'h18},
{8'h0D, 8'h25, 8'h5D},
{8'h1D, 8'h50, 8'hAE},
{8'h10, 8'h52, 8'hB9},
{8'h08, 8'h58, 8'hAE},
{8'h0F, 8'h4E, 8'hBB},
{8'h1D, 8'h4D, 8'hBA},
{8'h17, 8'h3C, 8'h8D},
{8'h03, 8'h20, 8'h6E},
{8'h18, 8'h40, 8'hA3},
{8'h20, 8'h54, 8'hB0},
{8'h0D, 8'h47, 8'h88},
{8'h05, 8'h06, 8'h2E},
{8'h03, 8'h00, 8'h14},
{8'h02, 8'h02, 8'h3E},
{8'h1E, 8'h3B, 8'h91},
{8'h17, 8'h56, 8'h8E},
{8'h30, 8'h6D, 8'h9D},
{8'h88, 8'hA3, 8'hC8},
{8'hE1, 8'hE6, 8'hDF},
{8'hF7, 8'hFF, 8'hFF},
{8'h8B, 8'hA2, 8'hC6},
{8'h22, 8'h4F, 8'hA3},
{8'h1C, 8'h3B, 8'h87},
{8'h04, 8'h01, 8'h25},
{8'h04, 8'h12, 8'h33},
{8'h00, 8'h14, 8'h37},
{8'h07, 8'h02, 8'h0A},
{8'h0A, 8'h02, 8'h2C},
{8'h02, 8'h00, 8'h0A},
{8'h8E, 8'h8F, 8'h73},
{8'hEB, 8'hEE, 8'hC2},
{8'hF0, 8'hF1, 8'hD0},
{8'hF5, 8'hF3, 8'hE4},
{8'hF3, 8'hF1, 8'hE3},
{8'hEE, 8'hEE, 8'hD7},
{8'hD4, 8'hD8, 8'hB1},
{8'hD6, 8'hD9, 8'hBB},
{8'hF4, 8'hF4, 8'hE4},
{8'hF8, 8'hF5, 8'hF0},
{8'hFA, 8'hF5, 8'hF1},
{8'hFB, 8'hF6, 8'hEB},
{8'hF7, 8'hF2, 8'hDD},
{8'hF4, 8'hEE, 8'hD0},
{8'hF8, 8'hEE, 8'hB8},
{8'hF3, 8'hEB, 8'hC9},
{8'hF3, 8'hEE, 8'hE5},
{8'hF8, 8'hF8, 8'hF9},
{8'hFC, 8'hFF, 8'hFC},
{8'hF9, 8'hFB, 8'hF4},
{8'hF9, 8'hF8, 8'hF1},
{8'hFE, 8'hFA, 8'hF7},
{8'hFA, 8'hFC, 8'hE1},
{8'hEE, 8'hF4, 8'hCF},
{8'hDE, 8'hE5, 8'hBB},
{8'hCD, 8'hD4, 8'hAA},
{8'hD3, 8'hD9, 8'hB8},
{8'h82, 8'h85, 8'h76},
{8'h77, 8'h77, 8'h7B},
{8'h7D, 8'h7B, 8'h89},
{8'h81, 8'h80, 8'h7E},
{8'h7B, 8'h7A, 8'h77},
{8'h7C, 8'h7B, 8'h79},
{8'h82, 8'h80, 8'h80},
{8'h81, 8'h7F, 8'h81},
{8'h7E, 8'h7C, 8'h7F},
{8'h81, 8'h7F, 8'h83},
{8'h7F, 8'h7D, 8'h82},
{8'h7E, 8'h7C, 8'h80},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'h7F, 8'h7D, 8'h7E},
{8'h82, 8'h80, 8'h81},
{8'h7C, 8'h7A, 8'h7B},
{8'h78, 8'h77, 8'h75},
{8'hA5, 8'hA5, 8'h9D},
{8'hFD, 8'hFD, 8'hEE},
{8'hFD, 8'hFE, 8'hE6},
{8'hED, 8'hEF, 8'hD2},
{8'hD8, 8'hD4, 8'hBF},
{8'hE6, 8'hE0, 8'hD1},
{8'hF0, 8'hEA, 8'hE2},
{8'hFD, 8'hFA, 8'hF5},
{8'hFE, 8'hFB, 8'hF4},
{8'hF9, 8'hF8, 8'hEA},
{8'hF1, 8'hF3, 8'hDB},
{8'hEE, 8'hF0, 8'hD2},
{8'hF0, 8'hEE, 8'hCB},
{8'hE9, 8'hE6, 8'hC5},
{8'hEB, 8'hE7, 8'hCC},
{8'hA9, 8'hA5, 8'h8E},
{8'hA9, 8'hA4, 8'h8D},
{8'hB5, 8'hB1, 8'h97},
{8'hC4, 8'hC1, 8'hA3},
{8'hD9, 8'hD7, 8'hB7},
{8'hC9, 8'hCA, 8'hB4},
{8'hBB, 8'hBD, 8'hA9},
{8'hD1, 8'hD2, 8'hC1},
{8'hDE, 8'hDE, 8'hD1},
{8'hF8, 8'hF8, 8'hED},
{8'hF3, 8'hF3, 8'hEB},
{8'hF0, 8'hEF, 8'hEB},
{8'hEE, 8'hED, 8'hE7},
{8'hE6, 8'hE3, 8'hCE},
{8'hF3, 8'hF0, 8'hE0},
{8'hFA, 8'hF6, 8'hF0},
{8'hFC, 8'hF7, 8'hF5},
{8'hFB, 8'hF7, 8'hF2},
{8'hFC, 8'hF9, 8'hE6},
{8'hFA, 8'hFA, 8'hD7},
{8'hED, 8'hF0, 8'hBE},
{8'hC6, 8'hCD, 8'h8D},
{8'h24, 8'h21, 8'h1D},
{8'h07, 8'h00, 8'h20},
{8'h05, 8'h03, 8'h1F},
{8'h00, 8'h04, 8'h21},
{8'h0D, 8'h25, 8'h64},
{8'h1D, 8'h51, 8'hB1},
{8'h11, 8'h52, 8'hBB},
{8'h15, 8'h52, 8'hBD},
{8'h27, 8'h55, 8'hAE},
{8'h17, 8'h33, 8'h78},
{8'h00, 8'h0B, 8'h49},
{8'h0D, 8'h34, 8'h7C},
{8'h1C, 8'h54, 8'hAC},
{8'h18, 8'h50, 8'hAF},
{8'h14, 8'h44, 8'hA3},
{8'h0A, 8'h18, 8'h49},
{8'h00, 8'h03, 8'h13},
{8'h00, 8'h02, 8'h24},
{8'h10, 8'h2B, 8'h70},
{8'h19, 8'h56, 8'hA5},
{8'h13, 8'h56, 8'hB9},
{8'h17, 8'h49, 8'hA7},
{8'h37, 8'h5B, 8'h8A},
{8'h6B, 8'h84, 8'hB1},
{8'h30, 8'h52, 8'h98},
{8'h1C, 8'h51, 8'hB3},
{8'h12, 8'h35, 8'h86},
{8'h01, 8'h00, 8'h26},
{8'h02, 8'h0F, 8'h3A},
{8'h08, 8'h20, 8'h55},
{8'h07, 8'h01, 8'h1F},
{8'h09, 8'h01, 8'h2B},
{8'h00, 8'h00, 8'h0A},
{8'h3A, 8'h3A, 8'h2D},
{8'hE5, 8'hE8, 8'hC7},
{8'hE5, 8'hE8, 8'hCE},
{8'hDA, 8'hDB, 8'hCC},
{8'hE0, 8'hE1, 8'hD2},
{8'hDE, 8'hE0, 8'hCA},
{8'hD7, 8'hDB, 8'hBA},
{8'hED, 8'hF0, 8'hD6},
{8'hF6, 8'hF4, 8'hE6},
{8'hF7, 8'hF5, 8'hED},
{8'hF8, 8'hF5, 8'hEA},
{8'hF7, 8'hF4, 8'hDE},
{8'hF5, 8'hF2, 8'hCF},
{8'hE6, 8'hE4, 8'hB5},
{8'hF0, 8'hEA, 8'h98},
{8'hF9, 8'hF3, 8'hB7},
{8'hFC, 8'hF8, 8'hDF},
{8'hFC, 8'hF9, 8'hF3},
{8'hFC, 8'hFC, 8'hF6},
{8'hFD, 8'hFD, 8'hF2},
{8'hF9, 8'hF8, 8'hE8},
{8'hEF, 8'hEC, 8'hDD},
{8'hED, 8'hEE, 8'hE3},
{8'hF8, 8'hFA, 8'hE9},
{8'hEB, 8'hEF, 8'hD5},
{8'hE6, 8'hEB, 8'hCD},
{8'hE1, 8'hE5, 8'hC8},
{8'h8E, 8'h92, 8'h7D},
{8'h79, 8'h7A, 8'h70},
{8'h7E, 8'h7E, 8'h7B},
{8'h74, 8'h73, 8'h70},
{8'h90, 8'h8F, 8'h8C},
{8'hA3, 8'hA2, 8'hA0},
{8'h7E, 8'h7C, 8'h7C},
{8'hBA, 8'hB8, 8'hBA},
{8'h82, 8'h80, 8'h83},
{8'h7E, 8'h7C, 8'h80},
{8'h81, 8'h7F, 8'h84},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'h8B, 8'h89, 8'h8A},
{8'h90, 8'h8E, 8'h8F},
{8'h7F, 8'h7D, 8'h7E},
{8'h82, 8'h81, 8'h80},
{8'hC6, 8'hC5, 8'hBE},
{8'hEE, 8'hEF, 8'hE1},
{8'hF6, 8'hF8, 8'hE3},
{8'hFB, 8'hFD, 8'hE2},
{8'hE9, 8'hE6, 8'hC7},
{8'hD6, 8'hD1, 8'hB8},
{8'hF1, 8'hEC, 8'hDD},
{8'hFB, 8'hF7, 8'hF0},
{8'hFA, 8'hF7, 8'hF1},
{8'hF7, 8'hF6, 8'hEC},
{8'hF5, 8'hF7, 8'hE7},
{8'hF5, 8'hF7, 8'hE2},
{8'hF5, 8'hF3, 8'hDB},
{8'hF0, 8'hEE, 8'hD5},
{8'hE9, 8'hE7, 8'hD0},
{8'hA9, 8'hA7, 8'h8F},
{8'h9F, 8'h9D, 8'h83},
{8'hB2, 8'hB1, 8'h91},
{8'hB1, 8'hB1, 8'h8D},
{8'hB2, 8'hB3, 8'h8E},
{8'h87, 8'h89, 8'h72},
{8'h8F, 8'h91, 8'h7D},
{8'hD2, 8'hD3, 8'hC1},
{8'hD1, 8'hD2, 8'hC2},
{8'hE3, 8'hE3, 8'hD6},
{8'hF0, 8'hF0, 8'hE5},
{8'hEB, 8'hEB, 8'hE2},
{8'hE0, 8'hDF, 8'hD6},
{8'hDB, 8'hD8, 8'hC9},
{8'hF3, 8'hF0, 8'hE4},
{8'hF7, 8'hF2, 8'hEB},
{8'hFC, 8'hF8, 8'hF2},
{8'hFE, 8'hFC, 8'hF0},
{8'hFE, 8'hFC, 8'hE3},
{8'hFB, 8'hFB, 8'hD6},
{8'hEF, 8'hF1, 8'hC0},
{8'h73, 8'h78, 8'h4F},
{8'h01, 8'h00, 8'h06},
{8'h07, 8'h02, 8'h26},
{8'h03, 8'h04, 8'h22},
{8'h00, 8'h05, 8'h2A},
{8'h0E, 8'h24, 8'h6B},
{8'h20, 8'h51, 8'hB2},
{8'h19, 8'h55, 8'hB9},
{8'h22, 8'h4C, 8'hB5},
{8'h14, 8'h2B, 8'h68},
{8'h00, 8'h03, 8'h28},
{8'h0F, 8'h1E, 8'h5C},
{8'h23, 8'h57, 8'hAB},
{8'h13, 8'h58, 8'hAD},
{8'h13, 8'h4F, 8'hAC},
{8'h1B, 8'h43, 8'hB0},
{8'h14, 8'h33, 8'h79},
{8'h00, 8'h0A, 8'h20},
{8'h00, 8'h02, 8'h0F},
{8'h0C, 8'h1D, 8'h50},
{8'h1C, 8'h51, 8'hB3},
{8'h09, 8'h4E, 8'hD6},
{8'h0C, 8'h52, 8'hD3},
{8'h13, 8'h54, 8'hAA},
{8'h1B, 8'h4A, 8'h9F},
{8'h1B, 8'h4E, 8'hAF},
{8'h11, 8'h52, 8'hBF},
{8'h0E, 8'h37, 8'h86},
{8'h00, 8'h00, 8'h21},
{8'h04, 8'h11, 8'h3C},
{8'h13, 8'h2D, 8'h6F},
{8'h04, 8'h00, 8'h2F},
{8'h08, 8'h01, 8'h2A},
{8'h04, 8'h01, 8'h17},
{8'h09, 8'h08, 8'h08},
{8'hAE, 8'hB0, 8'hA0},
{8'hE4, 8'hE6, 8'hD4},
{8'hD6, 8'hD7, 8'hC7},
{8'hDE, 8'hE0, 8'hCD},
{8'hEE, 8'hF0, 8'hDA},
{8'hD5, 8'hD9, 8'hC0},
{8'hE5, 8'hE8, 8'hD4},
{8'hF4, 8'hF5, 8'hE8},
{8'hF0, 8'hEE, 8'hE3},
{8'hF1, 8'hEF, 8'hDE},
{8'hF7, 8'hF7, 8'hD6},
{8'hFD, 8'hFD, 8'hCE},
{8'hE3, 8'hE5, 8'hA4},
{8'hD4, 8'hD3, 8'h62},
{8'hED, 8'hE9, 8'h95},
{8'hFD, 8'hF8, 8'hD0},
{8'hFC, 8'hF6, 8'hEA},
{8'hFA, 8'hF6, 8'hED},
{8'hF8, 8'hF6, 8'hE5},
{8'hF5, 8'hF4, 8'hDB},
{8'hF1, 8'hEF, 8'hD5},
{8'hE3, 8'hE4, 8'hDA},
{8'hF4, 8'hF6, 8'hEA},
{8'hFC, 8'hFE, 8'hEF},
{8'hF9, 8'hFC, 8'hE9},
{8'hEE, 8'hF1, 8'hDE},
{8'hB6, 8'hB9, 8'hA9},
{8'h8A, 8'h8B, 8'h81},
{8'h8E, 8'h8F, 8'h89},
{8'hB6, 8'hB5, 8'hB1},
{8'hCB, 8'hCA, 8'hC7},
{8'hEE, 8'hED, 8'hEB},
{8'hA2, 8'hA1, 8'hA0},
{8'hDE, 8'hDC, 8'hDE},
{8'h87, 8'h85, 8'h88},
{8'h7E, 8'h7C, 8'h80},
{8'h7E, 8'h7C, 8'h81},
{8'h7E, 8'h7C, 8'h7F},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'h7F, 8'h7E, 8'h7C},
{8'h7E, 8'h7C, 8'h7D},
{8'h7C, 8'h7A, 8'h7B},
{8'hA9, 8'hA8, 8'hA7},
{8'hEE, 8'hED, 8'hE8},
{8'hEF, 8'hEF, 8'hE3},
{8'hEC, 8'hED, 8'hDC},
{8'hF0, 8'hF2, 8'hD8},
{8'hEF, 8'hF1, 8'hB1},
{8'hD6, 8'hD6, 8'h9C},
{8'hDD, 8'hDC, 8'hB3},
{8'hE2, 8'hE0, 8'hC9},
{8'hEB, 8'hE9, 8'hDE},
{8'hF3, 8'hF1, 8'hED},
{8'hF2, 8'hF1, 8'hEE},
{8'hF2, 8'hF1, 8'hED},
{8'hF9, 8'hF7, 8'hEA},
{8'hF7, 8'hF4, 8'hE5},
{8'hEE, 8'hED, 8'hDB},
{8'hC9, 8'hC8, 8'hB1},
{8'h9E, 8'h9E, 8'h83},
{8'hB7, 8'hB7, 8'h98},
{8'hAF, 8'hAF, 8'h8D},
{8'h93, 8'h94, 8'h70},
{8'hAF, 8'hB0, 8'h9C},
{8'hE0, 8'hE1, 8'hD0},
{8'hCD, 8'hCE, 8'hBD},
{8'hA6, 8'hA7, 8'h97},
{8'hDA, 8'hDB, 8'hCD},
{8'hEA, 8'hEB, 8'hDE},
{8'hEA, 8'hEA, 8'hDE},
{8'hD3, 8'hD3, 8'hC7},
{8'hCA, 8'hC6, 8'hBE},
{8'hF4, 8'hF0, 8'hE8},
{8'hFA, 8'hF5, 8'hED},
{8'hF7, 8'hF4, 8'hE9},
{8'hF9, 8'hF6, 8'hE5},
{8'hF9, 8'hF8, 8'hDE},
{8'hFA, 8'hFA, 8'hD7},
{8'hD5, 8'hD7, 8'hAF},
{8'h1E, 8'h21, 8'h12},
{8'h03, 8'h00, 8'h12},
{8'h05, 8'h01, 8'h29},
{8'h01, 8'h01, 8'h21},
{8'h00, 8'h03, 8'h2A},
{8'h10, 8'h24, 8'h6E},
{8'h26, 8'h4D, 8'hAA},
{8'h17, 8'h48, 8'h9D},
{8'h0C, 8'h1C, 8'h67},
{8'h00, 8'h00, 8'h22},
{8'h06, 8'h0A, 8'h2C},
{8'h2A, 8'h41, 8'h98},
{8'h19, 8'h4F, 8'hC1},
{8'h0E, 8'h59, 8'hB6},
{8'h0F, 8'h4F, 8'hA1},
{8'h1A, 8'h44, 8'hA7},
{8'h20, 8'h43, 8'hA3},
{8'h02, 8'h0E, 8'h3D},
{8'h00, 8'h01, 8'h0B},
{8'h0A, 8'h16, 8'h3A},
{8'h21, 8'h47, 8'hAD},
{8'h0F, 8'h50, 8'hDB},
{8'h07, 8'h54, 8'hD1},
{8'h0B, 8'h59, 8'hB6},
{8'h15, 8'h54, 8'hB9},
{8'h10, 8'h50, 8'hBA},
{8'h0E, 8'h58, 8'hC3},
{8'h08, 8'h36, 8'h7B},
{8'h02, 8'h03, 8'h19},
{8'h03, 8'h14, 8'h39},
{8'h1D, 8'h3E, 8'h83},
{8'h07, 8'h08, 8'h40},
{8'h05, 8'h02, 8'h24},
{8'h09, 8'h06, 8'h22},
{8'h00, 8'h00, 8'h09},
{8'h5A, 8'h5A, 8'h5B},
{8'hEA, 8'hEB, 8'hE0},
{8'hE0, 8'hE2, 8'hCE},
{8'hE0, 8'hE5, 8'hCB},
{8'hF8, 8'hFC, 8'hE1},
{8'hE5, 8'hE9, 8'hD3},
{8'hD3, 8'hD7, 8'hC5},
{8'hD9, 8'hDA, 8'hCF},
{8'hE9, 8'hEA, 8'hDE},
{8'hE5, 8'hE5, 8'hD0},
{8'hE5, 8'hE7, 8'hC1},
{8'hF3, 8'hF7, 8'hC0},
{8'hD6, 8'hDB, 8'h92},
{8'hC2, 8'hC5, 8'h4A},
{8'hE1, 8'hE0, 8'h83},
{8'hFA, 8'hF5, 8'hC8},
{8'hFE, 8'hF7, 8'hE9},
{8'hFB, 8'hF4, 8'hEA},
{8'hFC, 8'hF9, 8'hE6},
{8'hF9, 8'hFA, 8'hDD},
{8'hF3, 8'hF5, 8'hD5},
{8'hCF, 8'hD3, 8'hB8},
{8'hE4, 8'hE8, 8'hD1},
{8'hFB, 8'hFD, 8'hEB},
{8'hF6, 8'hF7, 8'hEA},
{8'hF8, 8'hF8, 8'hF1},
{8'hFD, 8'hFD, 8'hFB},
{8'hF2, 8'hF1, 8'hF2},
{8'hEC, 8'hEB, 8'hEC},
{8'hFD, 8'hFC, 8'hF8},
{8'hF9, 8'hF8, 8'hF5},
{8'hF7, 8'hF6, 8'hF4},
{8'hF9, 8'hF8, 8'hF7},
{8'hC3, 8'hC1, 8'hC4},
{8'h7D, 8'h7B, 8'h7E},
{8'h7F, 8'h7D, 8'h81},
{8'h7E, 8'h7C, 8'h81},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'h7B, 8'h7A, 8'h77},
{8'h9E, 8'h9C, 8'h9C},
{8'hDD, 8'hDB, 8'hDC},
{8'hF6, 8'hF4, 8'hF5},
{8'hF4, 8'hF3, 8'hF0},
{8'hF3, 8'hF3, 8'hEA},
{8'hEC, 8'hED, 8'hDF},
{8'hE6, 8'hE8, 8'hCF},
{8'hCF, 8'hD5, 8'h7B},
{8'hD1, 8'hD6, 8'h83},
{8'hD7, 8'hD9, 8'h9D},
{8'hE6, 8'hE6, 8'hC3},
{8'hF4, 8'hF2, 8'hE2},
{8'hF1, 8'hEF, 8'hED},
{8'hF0, 8'hEE, 8'hF2},
{8'hD9, 8'hD6, 8'hDC},
{8'hC8, 8'hC5, 8'hC3},
{8'hF3, 8'hF0, 8'hEA},
{8'hFC, 8'hFA, 8'hEE},
{8'hED, 8'hEC, 8'hDA},
{8'hB7, 8'hB6, 8'h9F},
{8'h94, 8'h94, 8'h7A},
{8'hA3, 8'hA4, 8'h88},
{8'hE9, 8'hE9, 8'hD0},
{8'hFF, 8'hFF, 8'hF2},
{8'hCF, 8'hD0, 8'hC3},
{8'h8E, 8'h8F, 8'h82},
{8'hDC, 8'hDC, 8'hCF},
{8'hE6, 8'hE6, 8'hDB},
{8'hB7, 8'hB7, 8'hAB},
{8'hE2, 8'hE2, 8'hD7},
{8'hCF, 8'hCF, 8'hC4},
{8'h81, 8'h7C, 8'h78},
{8'h95, 8'h90, 8'h8B},
{8'hA9, 8'hA5, 8'h9B},
{8'hD7, 8'hD3, 8'hC6},
{8'hE5, 8'hE2, 8'hD0},
{8'hEF, 8'hEC, 8'hD7},
{8'hF6, 8'hF4, 8'hDC},
{8'h83, 8'h81, 8'h6D},
{8'h00, 8'h00, 8'h00},
{8'h01, 8'h00, 8'h1D},
{8'h01, 8'h00, 8'h28},
{8'h00, 8'h01, 8'h1E},
{8'h00, 8'h00, 8'h24},
{8'h1A, 8'h27, 8'h6C},
{8'h26, 8'h3F, 8'h8D},
{8'h01, 8'h15, 8'h4F},
{8'h00, 8'h05, 8'h29},
{8'h00, 8'h06, 8'h23},
{8'h17, 8'h2B, 8'h67},
{8'h28, 8'h4B, 8'hBE},
{8'h13, 8'h49, 8'hCE},
{8'h13, 8'h57, 8'hBE},
{8'h12, 8'h4F, 8'h9D},
{8'h16, 8'h48, 8'h9C},
{8'h22, 8'h49, 8'hBA},
{8'h0F, 8'h1E, 8'h6B},
{8'h00, 8'h00, 8'h18},
{8'h08, 8'h0D, 8'h2D},
{8'h29, 8'h46, 8'hA2},
{8'h19, 8'h52, 8'hCA},
{8'h09, 8'h52, 8'hB5},
{8'h0D, 8'h58, 8'hAC},
{8'h0D, 8'h52, 8'hB7},
{8'h10, 8'h54, 8'hBB},
{8'h0D, 8'h59, 8'hC0},
{8'h0D, 8'h3C, 8'h7D},
{8'h01, 8'h03, 8'h17},
{8'h03, 8'h17, 8'h3C},
{8'h21, 8'h4D, 8'h95},
{8'h0F, 8'h1A, 8'h57},
{8'h01, 8'h00, 8'h1A},
{8'h07, 8'h04, 8'h22},
{8'h01, 8'h00, 8'h1B},
{8'h13, 8'h12, 8'h20},
{8'hD5, 8'hD7, 8'hCF},
{8'hF1, 8'hF7, 8'hDC},
{8'hE3, 8'hEA, 8'hC6},
{8'hEB, 8'hF1, 8'hCE},
{8'hEC, 8'hF2, 8'hD7},
{8'hD9, 8'hDD, 8'hC9},
{8'hCE, 8'hD1, 8'hC4},
{8'hE1, 8'hE3, 8'hD7},
{8'hE4, 8'hE5, 8'hD3},
{8'hE3, 8'hE5, 8'hC3},
{8'hE0, 8'hE4, 8'hB0},
{8'hD4, 8'hD9, 8'h97},
{8'hD1, 8'hD7, 8'h6E},
{8'hE4, 8'hE5, 8'h97},
{8'hF3, 8'hEE, 8'hC8},
{8'hF5, 8'hEB, 8'hDE},
{8'hF1, 8'hEA, 8'hE0},
{8'hDF, 8'hDE, 8'hCA},
{8'hB8, 8'hBC, 8'hA2},
{8'hDF, 8'hE6, 8'hC9},
{8'hAC, 8'hB3, 8'h8A},
{8'hC8, 8'hCE, 8'hAB},
{8'hF1, 8'hF4, 8'hDE},
{8'hFB, 8'hFB, 8'hF3},
{8'hF7, 8'hF7, 8'hF8},
{8'hF7, 8'hF6, 8'hFC},
{8'hF9, 8'hF8, 8'hFF},
{8'hFA, 8'hF9, 8'hFD},
{8'hF5, 8'hF4, 8'hF0},
{8'hFA, 8'hF9, 8'hF6},
{8'hE9, 8'hE8, 8'hE6},
{8'hB5, 8'hB4, 8'hB4},
{8'h82, 8'h80, 8'h82},
{8'h79, 8'h77, 8'h7A},
{8'h82, 8'h80, 8'h84},
{8'h80, 8'h7E, 8'h83},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'h82, 8'h81, 8'h7D},
{8'hE6, 8'hE4, 8'hE3},
{8'hF4, 8'hF2, 8'hF3},
{8'hF2, 8'hF0, 8'hF1},
{8'hF7, 8'hF6, 8'hF4},
{8'hFB, 8'hFB, 8'hF5},
{8'hF6, 8'hF7, 8'hEB},
{8'hEE, 8'hF0, 8'hDC},
{8'hDA, 8'hDE, 8'h93},
{8'hCF, 8'hD1, 8'h8E},
{8'hE7, 8'hE8, 8'hB7},
{8'hF5, 8'hF4, 8'hD8},
{8'hF1, 8'hEF, 8'hE3},
{8'hEE, 8'hEC, 8'hE9},
{8'hB5, 8'hB3, 8'hB4},
{8'h87, 8'h85, 8'h87},
{8'h77, 8'h75, 8'h78},
{8'hA0, 8'h9F, 8'h9E},
{8'hE6, 8'hE5, 8'hDE},
{8'hF6, 8'hF6, 8'hE9},
{8'hD0, 8'hD1, 8'hC1},
{8'hC7, 8'hC8, 8'hB7},
{8'hF4, 8'hF4, 8'hE6},
{8'hFF, 8'hFF, 8'hF5},
{8'hD7, 8'hD7, 8'hD1},
{8'h7D, 8'h7D, 8'h76},
{8'hCE, 8'hCE, 8'hC7},
{8'hFF, 8'hFF, 8'hFB},
{8'hD6, 8'hD5, 8'hCE},
{8'h74, 8'h74, 8'h6B},
{8'hCF, 8'hD0, 8'hC6},
{8'hDE, 8'hDE, 8'hD6},
{8'h81, 8'h7C, 8'h7B},
{8'h7B, 8'h76, 8'h72},
{8'h99, 8'h95, 8'h8B},
{8'hE3, 8'hE0, 8'hD2},
{8'hF0, 8'hEC, 8'hDD},
{8'hF5, 8'hF1, 8'hE4},
{8'hEC, 8'hE7, 8'hDF},
{8'h33, 8'h2F, 8'h2D},
{8'h00, 8'h00, 8'h0B},
{8'h00, 8'h01, 8'h25},
{8'h01, 8'h00, 8'h25},
{8'h00, 8'h01, 8'h16},
{8'h03, 8'h04, 8'h23},
{8'h11, 8'h15, 8'h50},
{8'h06, 8'h09, 8'h42},
{8'h01, 8'h06, 8'h25},
{8'h02, 8'h05, 8'h18},
{8'h06, 8'h1B, 8'h4D},
{8'h19, 8'h4D, 8'hAA},
{8'h10, 8'h4F, 8'hC6},
{8'h14, 8'h4E, 8'hC5},
{8'h1C, 8'h50, 8'hB7},
{8'h13, 8'h4A, 8'hA2},
{8'h12, 8'h4E, 8'hA2},
{8'h1B, 8'h51, 8'hBD},
{8'h1E, 8'h3A, 8'h9B},
{8'h05, 8'h0A, 8'h37},
{8'h03, 8'h09, 8'h2E},
{8'h22, 8'h40, 8'h99},
{8'h1C, 8'h53, 8'hB9},
{8'h13, 8'h54, 8'hA8},
{8'h16, 8'h52, 8'hAF},
{8'h11, 8'h52, 8'hB3},
{8'h14, 8'h54, 8'hBA},
{8'h0F, 8'h54, 8'hC0},
{8'h18, 8'h40, 8'h8B},
{8'h02, 8'h04, 8'h25},
{8'h08, 8'h1F, 8'h51},
{8'h1B, 8'h54, 8'hA7},
{8'h15, 8'h2C, 8'h74},
{8'h03, 8'h01, 8'h15},
{8'h03, 8'h01, 8'h1C},
{8'h05, 8'h03, 8'h26},
{8'h02, 8'h01, 8'h17},
{8'h82, 8'h85, 8'h7D},
{8'hEF, 8'hF6, 8'hD2},
{8'hE4, 8'hEE, 8'hBE},
{8'hDF, 8'hE9, 8'hBB},
{8'hE9, 8'hF3, 8'hD1},
{8'hE8, 8'hEE, 8'hD4},
{8'hE4, 8'hE8, 8'hD8},
{8'hEE, 8'hF1, 8'hE6},
{8'hF3, 8'hF4, 8'hE7},
{8'hF1, 8'hF3, 8'hDB},
{8'hE3, 8'hE6, 8'hC0},
{8'hE7, 8'hEB, 8'hBA},
{8'hEB, 8'hF2, 8'hAF},
{8'hF5, 8'hF6, 8'hC7},
{8'hFB, 8'hF6, 8'hE1},
{8'hF8, 8'hF0, 8'hE8},
{8'hF3, 8'hEF, 8'hE3},
{8'hE9, 8'hEA, 8'hD9},
{8'h97, 8'hA0, 8'h8D},
{8'h95, 8'hA1, 8'h90},
{8'hA2, 8'hA9, 8'h86},
{8'hAB, 8'hAF, 8'h94},
{8'hE2, 8'hE4, 8'hD5},
{8'hF3, 8'hF4, 8'hEF},
{8'hFB, 8'hFB, 8'hFB},
{8'hFF, 8'hFF, 8'hFD},
{8'hFB, 8'hFC, 8'hF5},
{8'hF8, 8'hF9, 8'hEE},
{8'hF1, 8'hF0, 8'hEB},
{8'hD4, 8'hD3, 8'hD0},
{8'hA3, 8'hA2, 8'hA0},
{8'h78, 8'h76, 8'h76},
{8'h7B, 8'h79, 8'h7B},
{8'h80, 8'h7E, 8'h81},
{8'h7C, 8'h7A, 8'h7E},
{8'h7C, 8'h7A, 8'h7F},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'h7D, 8'h7C, 8'h77},
{8'h9C, 8'h9A, 8'h98},
{8'hA6, 8'hA4, 8'hA5},
{8'hA1, 8'h9F, 8'hA2},
{8'hA6, 8'hA5, 8'hA5},
{8'hD2, 8'hD1, 8'hCC},
{8'hF1, 8'hF1, 8'hE6},
{8'hF3, 8'hF3, 8'hE3},
{8'hED, 8'hEB, 8'hC8},
{8'hE6, 8'hE2, 8'hC5},
{8'hED, 8'hEA, 8'hD8},
{8'hDB, 8'hD7, 8'hCF},
{8'hEF, 8'hEB, 8'hE7},
{8'hDA, 8'hD8, 8'hD3},
{8'h81, 8'h81, 8'h76},
{8'h7E, 8'h7E, 8'h72},
{8'h83, 8'h80, 8'h87},
{8'h78, 8'h76, 8'h79},
{8'h82, 8'h81, 8'h7D},
{8'h88, 8'h88, 8'h7E},
{8'hB8, 8'hB8, 8'hAD},
{8'hFD, 8'hFD, 8'hF5},
{8'hFD, 8'hFC, 8'hF9},
{8'hDF, 8'hDD, 8'hDD},
{8'h84, 8'h82, 8'h82},
{8'hAF, 8'hAE, 8'hAD},
{8'hFF, 8'hFE, 8'hFC},
{8'hF9, 8'hF8, 8'hF5},
{8'h9B, 8'h9A, 8'h96},
{8'h7D, 8'h7D, 8'h78},
{8'hE5, 8'hE4, 8'hDF},
{8'hE0, 8'hDF, 8'hDA},
{8'h84, 8'h7E, 8'h7F},
{8'h7C, 8'h77, 8'h73},
{8'hC1, 8'hBD, 8'hB2},
{8'hF8, 8'hF5, 8'hE7},
{8'hF5, 8'hF0, 8'hE4},
{8'hFC, 8'hFA, 8'hF6},
{8'h9E, 8'h99, 8'h9C},
{8'h02, 8'h01, 8'h05},
{8'h01, 8'h03, 8'h1B},
{8'h00, 8'h00, 8'h29},
{8'h00, 8'h01, 8'h22},
{8'h01, 8'h02, 8'h10},
{8'h06, 8'h03, 8'h1A},
{8'h07, 8'h02, 8'h33},
{8'h05, 8'h00, 8'h2A},
{8'h05, 8'h03, 8'h0C},
{8'h0B, 8'h06, 8'h1A},
{8'h17, 8'h3A, 8'h8C},
{8'h08, 8'h57, 8'hCD},
{8'h01, 8'h5A, 8'hBF},
{8'h17, 8'h56, 8'hA9},
{8'h24, 8'h4A, 8'hAA},
{8'h15, 8'h42, 8'hAE},
{8'h0C, 8'h51, 8'hB5},
{8'h0E, 8'h58, 8'hB4},
{8'h1F, 8'h4C, 8'hB3},
{8'h11, 8'h23, 8'h63},
{8'h00, 8'h09, 8'h39},
{8'h15, 8'h3E, 8'h9A},
{8'h18, 8'h56, 8'hB7},
{8'h17, 8'h55, 8'hAC},
{8'h1C, 8'h4B, 8'hC1},
{8'h16, 8'h4F, 8'hB2},
{8'h1B, 8'h52, 8'hBC},
{8'h12, 8'h4E, 8'hC7},
{8'h23, 8'h42, 8'hA1},
{8'h04, 8'h04, 8'h38},
{8'h0C, 8'h29, 8'h70},
{8'h15, 8'h55, 8'hBA},
{8'h18, 8'h3E, 8'h92},
{8'h02, 8'h04, 8'h10},
{8'h04, 8'h04, 8'h1E},
{8'h01, 8'h00, 8'h2A},
{8'h01, 8'h01, 8'h1A},
{8'h22, 8'h27, 8'h20},
{8'hDC, 8'hE6, 8'hBA},
{8'hE8, 8'hF4, 8'hBB},
{8'hE1, 8'hED, 8'hB8},
{8'hE3, 8'hEF, 8'hC3},
{8'hE1, 8'hEB, 8'hCA},
{8'hE3, 8'hE8, 8'hD7},
{8'hF5, 8'hF7, 8'hF0},
{8'hF8, 8'hF9, 8'hF3},
{8'hFA, 8'hFB, 8'hEE},
{8'hF2, 8'hF3, 8'hDC},
{8'hE9, 8'hED, 8'hCE},
{8'hE8, 8'hEE, 8'hD1},
{8'hF0, 8'hF1, 8'hE1},
{8'hFB, 8'hF7, 8'hF4},
{8'hFE, 8'hFB, 8'hF8},
{8'hFC, 8'hFC, 8'hEF},
{8'hF8, 8'hFD, 8'hED},
{8'hCC, 8'hD9, 8'hCE},
{8'h83, 8'h92, 8'h8F},
{8'h8A, 8'h8E, 8'h81},
{8'h7E, 8'h80, 8'h78},
{8'h98, 8'h98, 8'h99},
{8'hF3, 8'hF2, 8'hF5},
{8'hF4, 8'hF5, 8'hF0},
{8'hFC, 8'hFE, 8'hEB},
{8'hEA, 8'hF1, 8'hC9},
{8'hEA, 8'hF1, 8'hC2},
{8'hDD, 8'hDC, 8'hD5},
{8'h84, 8'h82, 8'h80},
{8'h7A, 8'h79, 8'h78},
{8'h82, 8'h81, 8'h80},
{8'h83, 8'h81, 8'h83},
{8'h7B, 8'h79, 8'h7C},
{8'h80, 8'h7E, 8'h82},
{8'h83, 8'h81, 8'h86},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'h80, 8'h7F, 8'h7F},
{8'h7B, 8'h79, 8'h7A},
{8'h7B, 8'h79, 8'h7B},
{8'h7C, 8'h7A, 8'h7C},
{8'h7A, 8'h78, 8'h78},
{8'hD7, 8'hD6, 8'hD3},
{8'hF9, 8'hF8, 8'hF2},
{8'hF9, 8'hF8, 8'hF0},
{8'hFB, 8'hF8, 8'hF0},
{8'hF9, 8'hF5, 8'hF0},
{8'hE7, 8'hE3, 8'hE1},
{8'h89, 8'h86, 8'h87},
{8'hAE, 8'hAB, 8'hAC},
{8'hEC, 8'hEA, 8'hE8},
{8'hD2, 8'hD2, 8'hCC},
{8'h91, 8'h91, 8'h89},
{8'h7A, 8'h77, 8'h7D},
{8'h83, 8'h81, 8'h83},
{8'h7A, 8'h79, 8'h75},
{8'hA1, 8'hA1, 8'h97},
{8'hF8, 8'hF8, 8'hEF},
{8'hFE, 8'hFE, 8'hF8},
{8'hE1, 8'hDF, 8'hDF},
{8'h8C, 8'h8A, 8'h8E},
{8'h82, 8'h81, 8'h80},
{8'hEA, 8'hE9, 8'hE8},
{8'hFF, 8'hFF, 8'hFF},
{8'hD5, 8'hD3, 8'hD5},
{8'h7C, 8'h7A, 8'h7A},
{8'h85, 8'h84, 8'h82},
{8'hF0, 8'hEE, 8'hEB},
{8'hE8, 8'hE6, 8'hE2},
{8'h7F, 8'h7B, 8'h7B},
{8'h7E, 8'h7B, 8'h77},
{8'hE4, 8'hE2, 8'hDB},
{8'hFD, 8'hFC, 8'hF5},
{8'hFA, 8'hF7, 8'hF2},
{8'hEF, 8'hED, 8'hF2},
{8'h34, 8'h30, 8'h3E},
{8'h01, 8'h01, 8'h11},
{8'h02, 8'h03, 8'h22},
{8'h00, 8'h01, 8'h27},
{8'h00, 8'h01, 8'h22},
{8'h04, 8'h03, 8'h15},
{8'h0D, 8'h06, 8'h17},
{8'h0B, 8'h01, 8'h1F},
{8'h05, 8'h01, 8'h1E},
{8'h05, 8'h03, 8'h1B},
{8'h0D, 8'h24, 8'h62},
{8'h1D, 8'h52, 8'hB5},
{8'h0A, 8'h57, 8'hC9},
{8'h0B, 8'h5A, 8'hB9},
{8'h16, 8'h56, 8'hA7},
{8'h1F, 8'h4C, 8'hAB},
{8'h12, 8'h43, 8'hAF},
{8'h0F, 8'h50, 8'hB8},
{8'h0D, 8'h57, 8'hB7},
{8'h19, 8'h52, 8'hB9},
{8'h16, 8'h40, 8'h91},
{8'h01, 8'h13, 8'h57},
{8'h0C, 8'h39, 8'h91},
{8'h19, 8'h54, 8'hB0},
{8'h18, 8'h56, 8'hB4},
{8'h18, 8'h4F, 8'hC6},
{8'h12, 8'h50, 8'hB8},
{8'h1A, 8'h52, 8'hBB},
{8'h1A, 8'h4E, 8'hBB},
{8'h22, 8'h44, 8'hA2},
{8'h03, 8'h09, 8'h53},
{8'h11, 8'h38, 8'h8E},
{8'h15, 8'h56, 8'hC0},
{8'h16, 8'h4C, 8'hAC},
{8'h0C, 8'h10, 8'h25},
{8'h01, 8'h03, 8'h1C},
{8'h03, 8'h03, 8'h22},
{8'h04, 8'h03, 8'h19},
{8'h00, 8'h02, 8'h02},
{8'h8F, 8'h9E, 8'h85},
{8'hE4, 8'hFA, 8'hCB},
{8'hDE, 8'hF3, 8'hB9},
{8'hE2, 8'hF0, 8'hC4},
{8'hE0, 8'hED, 8'hC2},
{8'hE3, 8'hEE, 8'hC6},
{8'hEF, 8'hF7, 8'hD7},
{8'hF2, 8'hF7, 8'hE1},
{8'hE9, 8'hEE, 8'hD7},
{8'hEA, 8'hEE, 8'hD2},
{8'hEC, 8'hF2, 8'hD1},
{8'hE8, 8'hEB, 8'hDD},
{8'hED, 8'hEE, 8'hE7},
{8'hF0, 8'hEE, 8'hEC},
{8'hF9, 8'hF7, 8'hF4},
{8'hFB, 8'hFA, 8'hF5},
{8'hFC, 8'hFD, 8'hF7},
{8'hF1, 8'hF5, 8'hF5},
{8'h81, 8'h89, 8'h8E},
{8'h7C, 8'h7C, 8'h7E},
{8'h7C, 8'h7C, 8'h7E},
{8'h7C, 8'h7B, 8'h7D},
{8'hC0, 8'hC1, 8'hBE},
{8'hDE, 8'hE0, 8'hD5},
{8'hE9, 8'hED, 8'hD8},
{8'hE6, 8'hEB, 8'hCB},
{8'hD1, 8'hD7, 8'hB4},
{8'hAE, 8'hAE, 8'hA4},
{8'h7A, 8'h79, 8'h72},
{8'h80, 8'h7F, 8'h7A},
{8'h7E, 8'h7D, 8'h7A},
{8'h7F, 8'h7D, 8'h7E},
{8'hFF, 8'hD7, 8'h00},
{8'h7E, 8'h7C, 8'h81},
{8'h7F, 8'h7C, 8'h82},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'h7F, 8'h7D, 8'h82},
{8'h7F, 8'h7D, 8'h81},
{8'hFF, 8'hD7, 8'h00},
{8'h7C, 8'h7A, 8'h7C},
{8'h93, 8'h92, 8'h91},
{8'hF0, 8'hEF, 8'hED},
{8'hF6, 8'hF5, 8'hF2},
{8'hE8, 8'hE7, 8'hE4},
{8'hFA, 8'hFA, 8'hF6},
{8'hF3, 8'hF2, 8'hEF},
{8'hFB, 8'hFB, 8'hF9},
{8'hA5, 8'hA4, 8'hA3},
{8'h74, 8'h72, 8'h74},
{8'hAE, 8'hAC, 8'hAF},
{8'hB2, 8'hAF, 8'hB4},
{8'h7D, 8'h7B, 8'h81},
{8'h80, 8'h7E, 8'h82},
{8'h77, 8'h76, 8'h75},
{8'h91, 8'h90, 8'h8A},
{8'hEC, 8'hEC, 8'hE2},
{8'hFF, 8'hFF, 8'hF6},
{8'hD5, 8'hD5, 8'hCF},
{8'h88, 8'h86, 8'h86},
{8'h72, 8'h70, 8'h73},
{8'hAE, 8'hAE, 8'hA8},
{8'hFD, 8'hFC, 8'hF7},
{8'hF4, 8'hF3, 8'hF2},
{8'h97, 8'h95, 8'h98},
{8'h77, 8'h75, 8'h78},
{8'h8D, 8'h8C, 8'h8C},
{8'hFA, 8'hF9, 8'hF5},
{8'hEF, 8'hEE, 8'hE8},
{8'h86, 8'h82, 8'h81},
{8'h81, 8'h7F, 8'h7C},
{8'hE9, 8'hE8, 8'hE5},
{8'hFC, 8'hFB, 8'hFB},
{8'hFB, 8'hFC, 8'hFE},
{8'hAA, 8'hAA, 8'hB4},
{8'h03, 8'h03, 8'h14},
{8'h00, 8'h00, 8'h19},
{8'h04, 8'h00, 8'h21},
{8'h00, 8'h02, 8'h24},
{8'h00, 8'h03, 8'h23},
{8'h03, 8'h02, 8'h1B},
{8'h0B, 8'h02, 8'h13},
{8'h0B, 8'h01, 8'h16},
{8'h02, 8'h00, 8'h20},
{8'h04, 8'h0D, 8'h42},
{8'h07, 8'h44, 8'hAB},
{8'h16, 8'h58, 8'hBE},
{8'h12, 8'h51, 8'hB4},
{8'h16, 8'h52, 8'hB7},
{8'h14, 8'h51, 8'hB4},
{8'h14, 8'h51, 8'hB4},
{8'h0E, 8'h48, 8'hA9},
{8'h16, 8'h50, 8'hB1},
{8'h14, 8'h54, 8'hC3},
{8'h16, 8'h52, 8'hB9},
{8'h18, 8'h4E, 8'hAB},
{8'h05, 8'h29, 8'h7E},
{8'h11, 8'h32, 8'h83},
{8'h19, 8'h4E, 8'hA5},
{8'h19, 8'h56, 8'hB6},
{8'h11, 8'h55, 8'hBD},
{8'h0C, 8'h53, 8'hBD},
{8'h16, 8'h54, 8'hB8},
{8'h1F, 8'h51, 8'hAA},
{8'h1C, 8'h45, 8'h98},
{8'h03, 8'h18, 8'h6D},
{8'h16, 8'h47, 8'hA2},
{8'h16, 8'h55, 8'hB9},
{8'h13, 8'h55, 8'hBB},
{8'h13, 8'h19, 8'h44},
{8'h00, 8'h03, 8'h23},
{8'h00, 8'h02, 8'h1A},
{8'h04, 8'h01, 8'h15},
{8'h00, 8'h00, 8'h0A},
{8'h3F, 8'h48, 8'h4C},
{8'hDD, 8'hF0, 8'hD5},
{8'hE3, 8'hF6, 8'hC0},
{8'hDF, 8'hEE, 8'hC5},
{8'hE0, 8'hF1, 8'hBD},
{8'hE1, 8'hF2, 8'hB3},
{8'hE1, 8'hF0, 8'hB5},
{8'hE1, 8'hED, 8'hC1},
{8'hE6, 8'hEF, 8'hCE},
{8'hD4, 8'hDB, 8'hB9},
{8'hC7, 8'hCF, 8'hA8},
{8'hCF, 8'hCF, 8'hC1},
{8'hE4, 8'hE4, 8'hD9},
{8'hF3, 8'hF3, 8'hEA},
{8'hF3, 8'hF3, 8'hEE},
{8'hF9, 8'hF7, 8'hF8},
{8'hFE, 8'hFD, 8'hFF},
{8'hEE, 8'hEC, 8'hF0},
{8'h7E, 8'h7A, 8'h81},
{8'h7C, 8'h7C, 8'h7F},
{8'h7A, 8'h7A, 8'h79},
{8'h7F, 8'h80, 8'h7A},
{8'h8A, 8'h8C, 8'h81},
{8'hCF, 8'hD2, 8'hC5},
{8'hE2, 8'hE4, 8'hDA},
{8'hD6, 8'hD7, 8'hD2},
{8'h7B, 8'h7C, 8'h78},
{8'h95, 8'h95, 8'h89},
{8'h8E, 8'h8E, 8'h82},
{8'h7E, 8'h7E, 8'h75},
{8'h7F, 8'h7F, 8'h79},
{8'h7F, 8'h7E, 8'h7D},
{8'hFF, 8'hD7, 8'h00},
{8'h7F, 8'h7C, 8'h82},
{8'h7F, 8'h7C, 8'h83},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'h7F, 8'h7D, 8'h82},
{8'h7F, 8'h7D, 8'h81},
{8'hFF, 8'hD7, 8'h00},
{8'h79, 8'h77, 8'h79},
{8'hB3, 8'hB1, 8'hB1},
{8'hF6, 8'hF5, 8'hF3},
{8'hD8, 8'hD7, 8'hD4},
{8'h95, 8'h94, 8'h90},
{8'hEF, 8'hEF, 8'hEB},
{8'hF6, 8'hF5, 8'hF2},
{8'hFD, 8'hFD, 8'hFB},
{8'hCC, 8'hCB, 8'hCA},
{8'h7B, 8'h79, 8'h7B},
{8'h7D, 8'h7B, 8'h7E},
{8'h7E, 8'h7C, 8'h80},
{8'h7E, 8'h7C, 8'h81},
{8'h7D, 8'h7B, 8'h7E},
{8'h7D, 8'h7B, 8'h7B},
{8'hDA, 8'hD9, 8'hD4},
{8'hF4, 8'hF4, 8'hED},
{8'hB7, 8'hB6, 8'hAF},
{8'h83, 8'h82, 8'h7D},
{8'h79, 8'h78, 8'h77},
{8'h81, 8'h7F, 8'h81},
{8'hDB, 8'hDB, 8'hD5},
{8'hFE, 8'hFD, 8'hF9},
{8'hBC, 8'hBB, 8'hBB},
{8'h7C, 8'h7A, 8'h7D},
{8'hFF, 8'hD7, 8'h00},
{8'h96, 8'h95, 8'h94},
{8'hFB, 8'hFB, 8'hF6},
{8'hF6, 8'hF6, 8'hF0},
{8'h98, 8'h95, 8'h93},
{8'h79, 8'h77, 8'h75},
{8'hC8, 8'hC8, 8'hC5},
{8'hFF, 8'hFF, 8'hFF},
{8'hFE, 8'hFD, 8'hFE},
{8'h44, 8'h43, 8'h50},
{8'h01, 8'h00, 8'h14},
{8'h01, 8'h01, 8'h1A},
{8'h05, 8'h00, 8'h20},
{8'h01, 8'h01, 8'h23},
{8'h00, 8'h03, 8'h22},
{8'h02, 8'h02, 8'h1C},
{8'h04, 8'h01, 8'h17},
{8'h05, 8'h04, 8'h22},
{8'h00, 8'h02, 8'h31},
{8'h15, 8'h2F, 8'h6F},
{8'h19, 8'h57, 8'hBB},
{8'h17, 8'h56, 8'hBD},
{8'h11, 8'h51, 8'hB5},
{8'h17, 8'h55, 8'hB9},
{8'h14, 8'h51, 8'hB3},
{8'h15, 8'h51, 8'hB3},
{8'h0E, 8'h48, 8'hA9},
{8'h16, 8'h50, 8'hB2},
{8'h15, 8'h55, 8'hC3},
{8'h14, 8'h50, 8'hB7},
{8'h1C, 8'h52, 8'hAF},
{8'h17, 8'h46, 8'h9A},
{8'h09, 8'h2E, 8'h81},
{8'h1B, 8'h50, 8'hA9},
{8'h15, 8'h52, 8'hB3},
{8'h10, 8'h52, 8'hBA},
{8'h0D, 8'h53, 8'hBC},
{8'h16, 8'h54, 8'hB8},
{8'h1D, 8'h52, 8'hAD},
{8'h1B, 8'h43, 8'h98},
{8'h0A, 8'h28, 8'h7D},
{8'h1B, 8'h50, 8'hAC},
{8'h12, 8'h51, 8'hB5},
{8'h14, 8'h55, 8'hBC},
{8'h16, 8'h26, 8'h63},
{8'h00, 8'h00, 8'h2F},
{8'h00, 8'h01, 8'h25},
{8'h06, 8'h01, 8'h21},
{8'h0B, 8'h03, 8'h1A},
{8'h12, 8'h06, 8'h0D},
{8'h78, 8'h6E, 8'h58},
{8'hED, 8'hE9, 8'hBC},
{8'hE3, 8'hF1, 8'hC5},
{8'hE0, 8'hF1, 8'hBC},
{8'hE1, 8'hF2, 8'hB6},
{8'hE4, 8'hF2, 8'hBE},
{8'hD5, 8'hE0, 8'hBC},
{8'hA2, 8'hA9, 8'h93},
{8'h7F, 8'h84, 8'h70},
{8'h7B, 8'h80, 8'h67},
{8'h7C, 8'h7C, 8'h70},
{8'h9A, 8'h9A, 8'h91},
{8'hDF, 8'hDE, 8'hD8},
{8'hF9, 8'hF8, 8'hF4},
{8'hFC, 8'hFC, 8'hFB},
{8'hF9, 8'hF8, 8'hF9},
{8'hBA, 8'hB8, 8'hBD},
{8'h7D, 8'h7A, 8'h81},
{8'h7D, 8'h7C, 8'h80},
{8'h7B, 8'h7B, 8'h7A},
{8'h80, 8'h81, 8'h7B},
{8'hAE, 8'hB0, 8'hA6},
{8'hD7, 8'hD9, 8'hCE},
{8'hE6, 8'hE7, 8'hDE},
{8'hDB, 8'hDC, 8'hD6},
{8'h92, 8'h93, 8'h8E},
{8'h7A, 8'h7A, 8'h70},
{8'h94, 8'h94, 8'h8B},
{8'h88, 8'h87, 8'h81},
{8'h7D, 8'h7D, 8'h78},
{8'h7F, 8'h7D, 8'h7D},
{8'hFF, 8'hD7, 8'h00},
{8'h7F, 8'h7D, 8'h82},
{8'h7F, 8'h7C, 8'h83},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'h7F, 8'h7D, 8'h82},
{8'h7F, 8'h7D, 8'h81},
{8'h7E, 8'h7C, 8'h7F},
{8'h7D, 8'h7B, 8'h7D},
{8'hCD, 8'hCC, 8'hCB},
{8'hEC, 8'hEC, 8'hEA},
{8'h8F, 8'h8E, 8'h8B},
{8'h7A, 8'h79, 8'h74},
{8'hBC, 8'hBB, 8'hB7},
{8'hFB, 8'hFA, 8'hF7},
{8'hF5, 8'hF4, 8'hF2},
{8'hE1, 8'hE0, 8'hDF},
{8'h82, 8'h80, 8'h82},
{8'h7E, 8'h7C, 8'h7F},
{8'h80, 8'h7E, 8'h82},
{8'h7D, 8'h7B, 8'h80},
{8'h83, 8'h81, 8'h84},
{8'h85, 8'h83, 8'h84},
{8'hAF, 8'hAE, 8'hAC},
{8'h94, 8'h93, 8'h8F},
{8'h7B, 8'h7A, 8'h76},
{8'h7F, 8'h7D, 8'h7C},
{8'h81, 8'h7F, 8'h80},
{8'h95, 8'h93, 8'h95},
{8'hF5, 8'hF5, 8'hEF},
{8'hCD, 8'hCC, 8'hC8},
{8'h83, 8'h81, 8'h81},
{8'h7C, 8'h7A, 8'h7D},
{8'h7D, 8'h7B, 8'h7E},
{8'h99, 8'h98, 8'h97},
{8'hF9, 8'hF8, 8'hF3},
{8'hFA, 8'hFA, 8'hF4},
{8'hA1, 8'h9D, 8'h9D},
{8'h7A, 8'h77, 8'h77},
{8'h8C, 8'h8A, 8'h8A},
{8'hCD, 8'hCC, 8'hCD},
{8'h9F, 8'h9E, 8'hA5},
{8'h08, 8'h08, 8'h16},
{8'h04, 8'h04, 8'h18},
{8'h04, 8'h04, 8'h1E},
{8'h06, 8'h00, 8'h1D},
{8'h02, 8'h01, 8'h20},
{8'h00, 8'h03, 8'h21},
{8'h01, 8'h02, 8'h20},
{8'h03, 8'h04, 8'h21},
{8'h00, 8'h03, 8'h2D},
{8'h09, 8'h21, 8'h60},
{8'h1F, 8'h4E, 8'hA0},
{8'h14, 8'h53, 8'hB9},
{8'h13, 8'h53, 8'hB9},
{8'h14, 8'h54, 8'hB8},
{8'h14, 8'h53, 8'hB7},
{8'h13, 8'h50, 8'hB3},
{8'h15, 8'h51, 8'hB3},
{8'h0E, 8'h48, 8'hA9},
{8'h16, 8'h50, 8'hB2},
{8'h12, 8'h51, 8'hBE},
{8'h16, 8'h52, 8'hBA},
{8'h1B, 8'h52, 8'hB1},
{8'h1F, 8'h53, 8'hAB},
{8'h0E, 8'h3C, 8'h93},
{8'h18, 8'h4E, 8'hA9},
{8'h16, 8'h53, 8'hB5},
{8'h11, 8'h52, 8'hB9},
{8'h0E, 8'h52, 8'hBB},
{8'h16, 8'h54, 8'hB8},
{8'h1C, 8'h51, 8'hAF},
{8'h17, 8'h46, 8'h9D},
{8'h11, 8'h3A, 8'h92},
{8'h1C, 8'h52, 8'hB0},
{8'h16, 8'h54, 8'hB9},
{8'h11, 8'h52, 8'hBA},
{8'h1B, 8'h39, 8'h83},
{8'h00, 8'h01, 8'h34},
{8'h02, 8'h02, 8'h26},
{8'h08, 8'h01, 8'h25},
{8'h10, 8'h00, 8'h16},
{8'h37, 8'h11, 8'h10},
{8'h72, 8'h44, 8'h28},
{8'hB6, 8'h96, 8'h6A},
{8'hE6, 8'hF3, 8'hC4},
{8'hE0, 8'hF2, 8'hBA},
{8'hE1, 8'hF2, 8'hB6},
{8'hE6, 8'hF3, 8'hC3},
{8'hC6, 8'hCE, 8'hB4},
{8'h79, 8'h7D, 8'h74},
{8'h7C, 8'h7E, 8'h79},
{8'h7E, 8'h80, 8'h78},
{8'h82, 8'h81, 8'h7B},
{8'h7B, 8'h7B, 8'h75},
{8'h87, 8'h86, 8'h82},
{8'hBE, 8'hBD, 8'hBA},
{8'hCA, 8'hC9, 8'hC9},
{8'h98, 8'h96, 8'h99},
{8'h7F, 8'h7D, 8'h82},
{8'h7F, 8'h7D, 8'h82},
{8'h80, 8'h7F, 8'h83},
{8'h81, 8'h81, 8'h82},
{8'h7F, 8'h7F, 8'h7B},
{8'hB7, 8'hB8, 8'hB0},
{8'hED, 8'hEE, 8'hE5},
{8'hF9, 8'hF9, 8'hF4},
{8'hDE, 8'hDF, 8'hDA},
{8'h87, 8'h88, 8'h85},
{8'h7D, 8'h7D, 8'h76},
{8'h84, 8'h83, 8'h7E},
{8'h8F, 8'h8E, 8'h89},
{8'h7C, 8'h7B, 8'h78},
{8'h7E, 8'h7C, 8'h7D},
{8'hFF, 8'hD7, 8'h00},
{8'h7F, 8'h7D, 8'h82},
{8'h7F, 8'h7D, 8'h82},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'h7F, 8'h7D, 8'h82},
{8'h7F, 8'h7D, 8'h81},
{8'h7E, 8'h7C, 8'h7F},
{8'h82, 8'h7F, 8'h82},
{8'hB1, 8'hB0, 8'hAF},
{8'h97, 8'h96, 8'h94},
{8'h79, 8'h78, 8'h75},
{8'h81, 8'h80, 8'h7B},
{8'h84, 8'h83, 8'h7F},
{8'hDB, 8'hDA, 8'hD7},
{8'hFA, 8'hF9, 8'hF7},
{8'hEB, 8'hEA, 8'hE9},
{8'h89, 8'h87, 8'h89},
{8'h7B, 8'h79, 8'h7C},
{8'h7E, 8'h7C, 8'h80},
{8'h7F, 8'h7D, 8'h82},
{8'h81, 8'h7F, 8'h80},
{8'h7D, 8'h7B, 8'h7C},
{8'h76, 8'h74, 8'h75},
{8'h7C, 8'h7B, 8'h7B},
{8'h7D, 8'h7C, 8'h7C},
{8'h82, 8'h80, 8'h81},
{8'h7A, 8'h78, 8'h7A},
{8'hA5, 8'hA3, 8'hA4},
{8'hD1, 8'hD1, 8'hCB},
{8'h8A, 8'h89, 8'h85},
{8'h7D, 8'h7C, 8'h7B},
{8'h7D, 8'h7B, 8'h7E},
{8'h7C, 8'h7A, 8'h7D},
{8'h90, 8'h8F, 8'h8F},
{8'hF4, 8'hF4, 8'hF0},
{8'hF9, 8'hF9, 8'hF3},
{8'hA4, 8'hA0, 8'hA1},
{8'h77, 8'h74, 8'h75},
{8'h80, 8'h7E, 8'h7F},
{8'h80, 8'h7E, 8'h82},
{8'h2F, 8'h2F, 8'h36},
{8'h01, 8'h00, 8'h0F},
{8'h03, 8'h03, 8'h19},
{8'h04, 8'h03, 8'h1E},
{8'h06, 8'h00, 8'h1A},
{8'h04, 8'h01, 8'h1F},
{8'h00, 8'h02, 8'h21},
{8'h00, 8'h01, 8'h20},
{8'h02, 8'h03, 8'h26},
{8'h08, 8'h10, 8'h44},
{8'h1D, 8'h46, 8'h93},
{8'h18, 8'h54, 8'hB5},
{8'h0F, 8'h4F, 8'hB6},
{8'h12, 8'h51, 8'hB7},
{8'h15, 8'h55, 8'hB9},
{8'h13, 8'h51, 8'hB5},
{8'h14, 8'h51, 8'hB3},
{8'h14, 8'h50, 8'hB2},
{8'h10, 8'h4A, 8'hAC},
{8'h16, 8'h50, 8'hB2},
{8'h11, 8'h4F, 8'hBB},
{8'h16, 8'h52, 8'hBB},
{8'h18, 8'h52, 8'hB2},
{8'h1A, 8'h51, 8'hAC},
{8'h17, 8'h4F, 8'hA8},
{8'h0F, 8'h49, 8'hA6},
{8'h17, 8'h54, 8'hB5},
{8'h13, 8'h52, 8'hB9},
{8'h10, 8'h52, 8'hBA},
{8'h14, 8'h52, 8'hB7},
{8'h1A, 8'h51, 8'hB1},
{8'h16, 8'h48, 8'hA3},
{8'h14, 8'h47, 8'hA1},
{8'h19, 8'h50, 8'hAF},
{8'h17, 8'h55, 8'hBA},
{8'h10, 8'h53, 8'hBA},
{8'h19, 8'h43, 8'h90},
{8'h02, 8'h04, 8'h31},
{8'h04, 8'h02, 8'h1B},
{8'h06, 8'h01, 8'h1E},
{8'h22, 8'h09, 8'h19},
{8'h84, 8'h45, 8'h33},
{8'hA4, 8'h5A, 8'h2C},
{8'hAC, 8'h78, 8'h44},
{8'hE2, 8'hEE, 8'hBC},
{8'hE1, 8'hF4, 8'hBA},
{8'hE1, 8'hF2, 8'hB6},
{8'hE6, 8'hF3, 8'hC4},
{8'hB3, 8'hBB, 8'hA6},
{8'h79, 8'h7C, 8'h7C},
{8'h7C, 8'h7D, 8'h82},
{8'h7E, 8'h7F, 8'h81},
{8'h7D, 8'h7C, 8'h79},
{8'h7C, 8'h7B, 8'h78},
{8'h7C, 8'h7B, 8'h79},
{8'h7A, 8'h78, 8'h78},
{8'h80, 8'h7E, 8'h80},
{8'h7A, 8'h78, 8'h7B},
{8'h80, 8'h7E, 8'h81},
{8'h82, 8'h80, 8'h85},
{8'h7F, 8'h7E, 8'h83},
{8'h7F, 8'h7F, 8'h81},
{8'h7E, 8'h7F, 8'h7B},
{8'h73, 8'h75, 8'h6E},
{8'hAC, 8'hAD, 8'hA5},
{8'hF6, 8'hF7, 8'hF1},
{8'hB5, 8'hB6, 8'hB1},
{8'h76, 8'h76, 8'h75},
{8'h81, 8'h80, 8'h7D},
{8'h83, 8'h82, 8'h7F},
{8'h7F, 8'h7E, 8'h7C},
{8'h80, 8'h7E, 8'h7E},
{8'h7F, 8'h7D, 8'h7E},
{8'hFF, 8'hD7, 8'h00},
{8'h7F, 8'h7D, 8'h81},
{8'h7F, 8'h7D, 8'h82},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00}
};

    logic [23:0] Batt_rom [12511:0] = '{
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'h7C, 8'h7F, 8'h7F},
{8'h81, 8'h7C, 8'h81},
{8'h84, 8'h7A, 8'h83},
{8'h7F, 8'h7A, 8'h85},
{8'h74, 8'h7B, 8'h83},
{8'h76, 8'h7F, 8'h87},
{8'h7F, 8'h7E, 8'h88},
{8'h85, 8'h79, 8'h88},
{8'h7E, 8'h76, 8'h98},
{8'h81, 8'h7C, 8'h95},
{8'h7A, 8'h7A, 8'h85},
{8'h7B, 8'h7E, 8'h7B},
{8'h7A, 8'h7F, 8'h76},
{8'h81, 8'h84, 8'h7C},
{8'h80, 8'h7F, 8'h7D},
{8'h7C, 8'h7A, 8'h7B},
{8'h7F, 8'h7E, 8'h83},
{8'h7E, 8'h7D, 8'h82},
{8'h7E, 8'h7D, 8'h83},
{8'h80, 8'h7F, 8'h85},
{8'h7E, 8'h7D, 8'h83},
{8'h7E, 8'h7D, 8'h82},
{8'h7E, 8'h7D, 8'h82},
{8'h7E, 8'h7D, 8'h83},
{8'h86, 8'h80, 8'h88},
{8'h81, 8'h7C, 8'h84},
{8'h7D, 8'h7A, 8'h81},
{8'h7E, 8'h7D, 8'h82},
{8'h7B, 8'h7D, 8'h80},
{8'h7D, 8'h81, 8'h82},
{8'h7C, 8'h83, 8'h81},
{8'h79, 8'h80, 8'h7F},
{8'h7D, 8'h79, 8'h8D},
{8'h7E, 8'h7B, 8'h88},
{8'h7E, 8'h7E, 8'h7F},
{8'h7F, 8'h80, 8'h77},
{8'h7E, 8'h80, 8'h74},
{8'h7E, 8'h7F, 8'h79},
{8'h7E, 8'h7D, 8'h82},
{8'h7F, 8'h7D, 8'h86},
{8'h82, 8'h83, 8'h70},
{8'h7E, 8'h7E, 8'h77},
{8'h78, 8'h76, 8'h7E},
{8'h7C, 8'h78, 8'h84},
{8'h7E, 8'h7B, 8'h80},
{8'h7C, 8'h7A, 8'h79},
{8'h7F, 8'h7D, 8'h82},
{8'h80, 8'h7D, 8'h88},
{8'h81, 8'h80, 8'h79},
{8'h96, 8'h95, 8'h8F},
{8'h7C, 8'h7B, 8'h7B},
{8'h7E, 8'h7C, 8'h82},
{8'h7F, 8'h7C, 8'h82},
{8'h7F, 8'h7D, 8'h7F},
{8'h7F, 8'h7E, 8'h79},
{8'h7F, 8'h7F, 8'h78},
{8'h7F, 8'h7D, 8'h7F},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'h7E, 8'h7D, 8'h80},
{8'h7A, 8'h80, 8'h82},
{8'h80, 8'h7C, 8'h82},
{8'h84, 8'h7A, 8'h83},
{8'h82, 8'h7C, 8'h83},
{8'h7A, 8'h7E, 8'h81},
{8'h79, 8'h7F, 8'h7F},
{8'h7F, 8'h7D, 8'h7E},
{8'h86, 8'h79, 8'h7D},
{8'h7F, 8'h7B, 8'h7E},
{8'h81, 8'h7F, 8'h81},
{8'h7D, 8'h7C, 8'h7C},
{8'h7E, 8'h7F, 8'h7C},
{8'h7D, 8'h7D, 8'h7D},
{8'h81, 8'h7F, 8'h84},
{8'h7E, 8'h7C, 8'h85},
{8'h7E, 8'h7A, 8'h86},
{8'h80, 8'h7E, 8'h7D},
{8'h7F, 8'h7D, 8'h7B},
{8'h7D, 8'h7B, 8'h79},
{8'h7C, 8'h7A, 8'h78},
{8'h7A, 8'h77, 8'h75},
{8'h79, 8'h77, 8'h75},
{8'h79, 8'h77, 8'h75},
{8'h7A, 8'h77, 8'h75},
{8'h80, 8'h79, 8'h78},
{8'h81, 8'h7A, 8'h79},
{8'h80, 8'h7B, 8'h7A},
{8'h80, 8'h7D, 8'h7C},
{8'h80, 8'h7E, 8'h7D},
{8'h7E, 8'h7F, 8'h7D},
{8'h7F, 8'h82, 8'h7D},
{8'h7B, 8'h7E, 8'h7B},
{8'h7E, 8'h79, 8'h84},
{8'h7F, 8'h7A, 8'h83},
{8'h7F, 8'h7C, 8'h80},
{8'h7F, 8'h7E, 8'h7C},
{8'h7F, 8'h7E, 8'h7B},
{8'h7F, 8'h7E, 8'h7E},
{8'h7E, 8'h7E, 8'h81},
{8'h7E, 8'h7D, 8'h81},
{8'h7F, 8'h7F, 8'h73},
{8'h87, 8'h86, 8'h82},
{8'h96, 8'h94, 8'h97},
{8'h89, 8'h88, 8'h87},
{8'h85, 8'h85, 8'h7A},
{8'h7B, 8'h7C, 8'h6E},
{8'h7A, 8'h79, 8'h74},
{8'h7D, 8'h7B, 8'h7F},
{8'h85, 8'h85, 8'h7E},
{8'h9B, 8'h9A, 8'h96},
{8'h7B, 8'h79, 8'h7B},
{8'h7E, 8'h7C, 8'h82},
{8'h7F, 8'h7C, 8'h83},
{8'h7F, 8'h7D, 8'h81},
{8'h7F, 8'h7E, 8'h7C},
{8'h7F, 8'h7E, 8'h7A},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'h7E, 8'h7D, 8'h81},
{8'h77, 8'h80, 8'h87},
{8'h7E, 8'h7D, 8'h85},
{8'h84, 8'h7A, 8'h81},
{8'h84, 8'h7B, 8'h7D},
{8'h81, 8'h82, 8'h7B},
{8'h75, 8'h78, 8'h6D},
{8'h79, 8'h74, 8'h67},
{8'h86, 8'h78, 8'h6B},
{8'h83, 8'h81, 8'h67},
{8'h83, 8'h83, 8'h6C},
{8'h7C, 8'h79, 8'h6D},
{8'h7E, 8'h7A, 8'h79},
{8'h85, 8'h7F, 8'h87},
{8'h80, 8'h79, 8'h86},
{8'h7F, 8'h78, 8'h87},
{8'h7C, 8'h76, 8'h82},
{8'h7A, 8'h76, 8'h68},
{8'h7C, 8'h78, 8'h67},
{8'h8C, 8'h88, 8'h78},
{8'hA3, 8'h9E, 8'h8E},
{8'hB2, 8'hAE, 8'h9E},
{8'hB2, 8'hAE, 8'h9E},
{8'hB2, 8'hAE, 8'h9E},
{8'hB2, 8'hAE, 8'h9E},
{8'hA8, 8'hA1, 8'h90},
{8'h93, 8'h8C, 8'h7C},
{8'h86, 8'h7E, 8'h70},
{8'h85, 8'h7E, 8'h72},
{8'h7E, 8'h77, 8'h6E},
{8'h7E, 8'h79, 8'h71},
{8'h7E, 8'h7A, 8'h73},
{8'h81, 8'h7E, 8'h79},
{8'h7F, 8'h79, 8'h74},
{8'h80, 8'h79, 8'h77},
{8'h81, 8'h7A, 8'h7F},
{8'h80, 8'h7B, 8'h82},
{8'h80, 8'h7C, 8'h85},
{8'h7F, 8'h7C, 8'h83},
{8'h7E, 8'h7E, 8'h80},
{8'h7D, 8'h7D, 8'h7B},
{8'h83, 8'h82, 8'h7F},
{8'hB6, 8'hB4, 8'hB4},
{8'hBE, 8'hBD, 8'hB9},
{8'hD2, 8'hD4, 8'hC2},
{8'hE8, 8'hEB, 8'hCB},
{8'hC9, 8'hCD, 8'hAA},
{8'h93, 8'h95, 8'h7F},
{8'h7D, 8'h7D, 8'h75},
{8'h89, 8'h88, 8'h82},
{8'hA3, 8'hA2, 8'h9E},
{8'h7A, 8'h78, 8'h79},
{8'h80, 8'h7D, 8'h82},
{8'h7F, 8'h7C, 8'h83},
{8'h7F, 8'h7D, 8'h81},
{8'hFF, 8'hD7, 8'h00},
{8'h7F, 8'h7D, 8'h7D},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'h7E, 8'h7D, 8'h81},
{8'h76, 8'h80, 8'h88},
{8'h7D, 8'h7D, 8'h84},
{8'h86, 8'h7A, 8'h7D},
{8'h85, 8'h79, 8'h73},
{8'h7E, 8'h7B, 8'h6B},
{8'hA2, 8'hA3, 8'h8D},
{8'hD0, 8'hCA, 8'hB3},
{8'hE7, 8'hDD, 8'hC7},
{8'hE0, 8'hDF, 8'hC0},
{8'hD2, 8'hD0, 8'hB7},
{8'hC2, 8'hBB, 8'hB0},
{8'hA5, 8'h9A, 8'h9A},
{8'h82, 8'h75, 8'h7B},
{8'h84, 8'h79, 8'h7D},
{8'h79, 8'h73, 8'h71},
{8'h99, 8'h96, 8'h8D},
{8'hC3, 8'hBD, 8'hA3},
{8'hE4, 8'hDF, 8'hC3},
{8'hFA, 8'hF7, 8'hDC},
{8'hFF, 8'hFD, 8'hE1},
{8'hFF, 8'hFF, 8'hE3},
{8'hFF, 8'hFE, 8'hE2},
{8'hFF, 8'hFE, 8'hE3},
{8'hFF, 8'hFD, 8'hE1},
{8'hF9, 8'hF3, 8'hD2},
{8'hF4, 8'hF0, 8'hD1},
{8'hF0, 8'hEC, 8'hD0},
{8'hDB, 8'hD7, 8'hBF},
{8'hBB, 8'hB4, 8'hA0},
{8'h98, 8'h8E, 8'h7E},
{8'h98, 8'h8D, 8'h81},
{8'h95, 8'h8B, 8'h80},
{8'h8C, 8'h84, 8'h6E},
{8'h87, 8'h7E, 8'h71},
{8'h82, 8'h79, 8'h79},
{8'h82, 8'h79, 8'h85},
{8'h81, 8'h79, 8'h88},
{8'h81, 8'h7D, 8'h87},
{8'h7F, 8'h7D, 8'h7F},
{8'h7E, 8'h7E, 8'h7A},
{8'h80, 8'h7E, 8'h83},
{8'h81, 8'h7F, 8'h82},
{8'h7C, 8'h7B, 8'h73},
{8'h8D, 8'h90, 8'h73},
{8'hE6, 8'hEC, 8'hBC},
{8'hF5, 8'hFC, 8'hC8},
{8'hF0, 8'hF5, 8'hCF},
{8'h9C, 8'h9E, 8'h89},
{8'h87, 8'h87, 8'h7C},
{8'hA3, 8'hA3, 8'h9B},
{8'h77, 8'h77, 8'h71},
{8'h7F, 8'h7E, 8'h7B},
{8'h7E, 8'h7C, 8'h7C},
{8'h7E, 8'h7D, 8'h7D},
{8'h7E, 8'h7C, 8'h7E},
{8'h7F, 8'h7D, 8'h7F},
{8'h7E, 8'h7C, 8'h7F},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'h7E, 8'h7C, 8'h7F},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'h7E, 8'h7D, 8'h80},
{8'h7A, 8'h83, 8'h88},
{8'h83, 8'h80, 8'h83},
{8'h8A, 8'h78, 8'h77},
{8'h81, 8'h70, 8'h65},
{8'hC3, 8'hBC, 8'hA7},
{8'hFA, 8'hF9, 8'hE1},
{8'hD3, 8'hCE, 8'hB7},
{8'hB2, 8'hA7, 8'h95},
{8'h9D, 8'h98, 8'h8B},
{8'h9C, 8'h93, 8'h8B},
{8'hAF, 8'hA1, 8'h9C},
{8'hB9, 8'hA7, 8'hA2},
{8'hA4, 8'h93, 8'h8A},
{8'h9C, 8'h90, 8'h7D},
{8'hD3, 8'hD0, 8'hB2},
{8'hF9, 8'hF8, 8'hD3},
{8'hFF, 8'hFF, 8'hDC},
{8'hFF, 8'hFE, 8'hDB},
{8'hF0, 8'hEB, 8'hC7},
{8'hEF, 8'hEB, 8'hC7},
{8'hF7, 8'hF3, 8'hCF},
{8'hFF, 8'hFC, 8'hD9},
{8'hFF, 8'hFF, 8'hDC},
{8'hFF, 8'hFC, 8'hD7},
{8'hF5, 8'hEF, 8'hC5},
{8'hEB, 8'hE3, 8'hBA},
{8'hF3, 8'hED, 8'hC8},
{8'hFE, 8'hF9, 8'hD8},
{8'hFF, 8'hFF, 8'hE3},
{8'hFC, 8'hF5, 8'hDD},
{8'hE6, 8'hD9, 8'hC5},
{8'hDC, 8'hCD, 8'hB9},
{8'hF1, 8'hE8, 8'hC5},
{8'hDD, 8'hD3, 8'hB9},
{8'h7E, 8'h71, 8'h68},
{8'h81, 8'h76, 8'h7B},
{8'h83, 8'h7A, 8'h85},
{8'h81, 8'h7B, 8'h83},
{8'h7C, 8'h7A, 8'h7B},
{8'h81, 8'h81, 8'h7E},
{8'h7E, 8'h7C, 8'h82},
{8'h7C, 8'h7A, 8'h80},
{8'h7E, 8'h7D, 8'h78},
{8'h99, 8'h9B, 8'h81},
{8'hF0, 8'hF5, 8'hC4},
{8'hEF, 8'hF7, 8'hBD},
{8'hF2, 8'hF8, 8'hC8},
{8'hBC, 8'hC0, 8'h9C},
{8'hAC, 8'hAD, 8'h99},
{8'hB8, 8'hBA, 8'hA7},
{8'h82, 8'h84, 8'h71},
{8'h7C, 8'h7D, 8'h6C},
{8'h86, 8'h87, 8'h7A},
{8'h80, 8'h80, 8'h76},
{8'h80, 8'h7F, 8'h79},
{8'h78, 8'h77, 8'h74},
{8'h7F, 8'h7D, 8'h7F},
{8'hFF, 8'hD7, 8'h00},
{8'h7D, 8'h7B, 8'h7E},
{8'h7C, 8'h7A, 8'h7D},
{8'h7E, 8'h7C, 8'h7F},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'h7D, 8'h7C, 8'h7F},
{8'h7E, 8'h82, 8'h80},
{8'h86, 8'h7D, 8'h78},
{8'h81, 8'h68, 8'h61},
{8'hB8, 8'hA4, 8'h96},
{8'hEA, 8'hE4, 8'hCF},
{8'h9B, 8'h99, 8'h85},
{8'h7A, 8'h77, 8'h67},
{8'h7F, 8'h76, 8'h6E},
{8'h83, 8'h7A, 8'h81},
{8'h84, 8'h77, 8'h7A},
{8'h85, 8'h72, 8'h6C},
{8'h82, 8'h6C, 8'h5B},
{8'hBC, 8'hAB, 8'h8E},
{8'hEC, 8'hE2, 8'hBA},
{8'hF0, 8'hEC, 8'hBC},
{8'hF8, 8'hF9, 8'hC8},
{8'hFC, 8'hF9, 8'hD3},
{8'hFF, 8'hFD, 8'hD9},
{8'hF9, 8'hF6, 8'hD1},
{8'hF0, 8'hED, 8'hC7},
{8'hEA, 8'hE4, 8'hBE},
{8'hFC, 8'hF9, 8'hD3},
{8'hFF, 8'hFE, 8'hD7},
{8'hFE, 8'hFD, 8'hD6},
{8'hFD, 8'hFB, 8'hCF},
{8'hFE, 8'hFC, 8'hD1},
{8'hFB, 8'hF9, 8'hCF},
{8'hF5, 8'hEF, 8'hC8},
{8'hEE, 8'hE6, 8'hC2},
{8'hF8, 8'hEF, 8'hCF},
{8'hFF, 8'hFC, 8'hDD},
{8'hF5, 8'hE9, 8'hCA},
{8'hE9, 8'hDC, 8'hB2},
{8'hEF, 8'hE5, 8'hC0},
{8'h92, 8'h84, 8'h6B},
{8'h82, 8'h77, 8'h68},
{8'h84, 8'h7B, 8'h77},
{8'h85, 8'h80, 8'h80},
{8'h82, 8'h7F, 8'h81},
{8'h7F, 8'h7E, 8'h7F},
{8'h80, 8'h7F, 8'h81},
{8'h7B, 8'h78, 8'h7F},
{8'h79, 8'h77, 8'h7C},
{8'hAD, 8'hAE, 8'hA1},
{8'hC5, 8'hC9, 8'hA5},
{8'hE9, 8'hF1, 8'hBD},
{8'hEE, 8'hF6, 8'hC1},
{8'hED, 8'hF3, 8'hC4},
{8'hEF, 8'hF3, 8'hCF},
{8'hF2, 8'hF6, 8'hD2},
{8'hE2, 8'hE5, 8'hC1},
{8'hD0, 8'hD4, 8'hB1},
{8'hDF, 8'hE2, 8'hC3},
{8'hD7, 8'hD9, 8'hC1},
{8'hD1, 8'hD3, 8'hC1},
{8'hAA, 8'hAB, 8'h9F},
{8'h7D, 8'h7B, 8'h7D},
{8'hFF, 8'hD7, 8'h00},
{8'h7E, 8'h7C, 8'h7F},
{8'h81, 8'h7F, 8'h82},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'h7B, 8'h79, 8'h6F},
{8'h83, 8'h73, 8'h68},
{8'h93, 8'h76, 8'h68},
{8'hDD, 8'hC5, 8'hB4},
{8'h92, 8'h84, 8'h72},
{8'h7D, 8'h7C, 8'h6E},
{8'h7D, 8'h7D, 8'h79},
{8'h82, 8'h7E, 8'h84},
{8'h80, 8'h76, 8'h81},
{8'h88, 8'h7B, 8'h7A},
{8'h84, 8'h71, 8'h5E},
{8'hBB, 8'hA3, 8'h7F},
{8'hFF, 8'hF6, 8'hC7},
{8'hF3, 8'hE9, 8'hB8},
{8'hE9, 8'hE4, 8'hB9},
{8'hF6, 8'hF4, 8'hCF},
{8'hF6, 8'hF4, 8'hCF},
{8'hFD, 8'hFD, 8'hD9},
{8'hFF, 8'hFF, 8'hDA},
{8'hFE, 8'hFC, 8'hD7},
{8'hFC, 8'hFA, 8'hD6},
{8'hFB, 8'hF8, 8'hD2},
{8'hFF, 8'hFE, 8'hD9},
{8'hFF, 8'hFF, 8'hD9},
{8'hF9, 8'hF8, 8'hCD},
{8'hF9, 8'hF8, 8'hCF},
{8'hF9, 8'hF7, 8'hCD},
{8'hF5, 8'hF3, 8'hC9},
{8'hF4, 8'hF0, 8'hC7},
{8'hDD, 8'hD2, 8'hAA},
{8'hE9, 8'hDD, 8'hB5},
{8'hF7, 8'hEF, 8'hC8},
{8'hFC, 8'hF1, 8'hC5},
{8'hE2, 8'hD2, 8'hA6},
{8'h9B, 8'h8D, 8'h64},
{8'hB0, 8'hA7, 8'h84},
{8'h86, 8'h7F, 8'h67},
{8'h81, 8'h7B, 8'h72},
{8'h7E, 8'h7B, 8'h7D},
{8'h7E, 8'h7C, 8'h85},
{8'h80, 8'h7F, 8'h7B},
{8'h85, 8'h83, 8'h89},
{8'h7C, 8'h78, 8'h89},
{8'h81, 8'h7E, 8'h85},
{8'h81, 8'h82, 8'h71},
{8'hE3, 8'hE8, 8'hC1},
{8'hEE, 8'hF5, 8'hC2},
{8'hEC, 8'hF3, 8'hBE},
{8'hF1, 8'hF8, 8'hC5},
{8'hEE, 8'hF4, 8'hC0},
{8'hEE, 8'hF6, 8'hBF},
{8'hF1, 8'hF9, 8'hC2},
{8'hF2, 8'hF8, 8'hC9},
{8'hF6, 8'hFA, 8'hD3},
{8'hD2, 8'hD5, 8'hB6},
{8'hD7, 8'hD9, 8'hC2},
{8'hAC, 8'hAA, 8'hAC},
{8'h7A, 8'h78, 8'h7B},
{8'h81, 8'h7F, 8'h82},
{8'h81, 8'h7F, 8'h82},
{8'h80, 8'h7E, 8'h81},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'h7F, 8'h7D, 8'h7F},
{8'h7F, 8'h7D, 8'h7F},
{8'hFF, 8'hD7, 8'h00},
{8'h7F, 8'h7D, 8'h81},
{8'h7F, 8'h7D, 8'h81},
{8'hFF, 8'hD7, 8'h00},
{8'h7F, 8'h7D, 8'h7F},
{8'h7F, 8'h7D, 8'h7E},
{8'h86, 8'h80, 8'h70},
{8'h85, 8'h6C, 8'h5C},
{8'hB0, 8'h8F, 8'h7E},
{8'hA4, 8'h89, 8'h77},
{8'h84, 8'h76, 8'h66},
{8'h7E, 8'h7C, 8'h76},
{8'h79, 8'h7C, 8'h84},
{8'h7E, 8'h7F, 8'h8C},
{8'h82, 8'h7A, 8'h7D},
{8'h8B, 8'h75, 8'h6A},
{8'h98, 8'h7E, 8'h5E},
{8'hDD, 8'hCD, 8'h9B},
{8'hFE, 8'hF6, 8'hC1},
{8'hF2, 8'hE4, 8'hB7},
{8'hFF, 8'hFB, 8'hDB},
{8'hF2, 8'hEF, 8'hD6},
{8'hF2, 8'hF2, 8'hCF},
{8'hF6, 8'hF5, 8'hD0},
{8'hF9, 8'hF9, 8'hD3},
{8'hFC, 8'hFC, 8'hD7},
{8'hFD, 8'hFD, 8'hD9},
{8'hFF, 8'hFF, 8'hDC},
{8'hFE, 8'hFE, 8'hD9},
{8'hFF, 8'hFF, 8'hD9},
{8'hFD, 8'hFD, 8'hD9},
{8'hEC, 8'hEA, 8'hC3},
{8'hF2, 8'hEF, 8'hC6},
{8'hF5, 8'hF2, 8'hCA},
{8'hEF, 8'hE8, 8'hBE},
{8'hF8, 8'hF1, 8'hC6},
{8'hF1, 8'hE7, 8'hBC},
{8'hEF, 8'hE6, 8'hB9},
{8'hF1, 8'hDF, 8'hB2},
{8'hFA, 8'hEB, 8'hBB},
{8'hC6, 8'hB9, 8'h87},
{8'hF1, 8'hE9, 8'hB9},
{8'hD9, 8'hD3, 8'hAF},
{8'h7F, 8'h79, 8'h66},
{8'h7C, 8'h78, 8'h77},
{8'h7B, 8'h79, 8'h80},
{8'h79, 8'h79, 8'h6D},
{8'h7D, 8'h7B, 8'h7E},
{8'h7D, 8'h78, 8'h8D},
{8'h7D, 8'h79, 8'h8A},
{8'h89, 8'h88, 8'h84},
{8'hDA, 8'hDD, 8'hBE},
{8'hED, 8'hF3, 8'hC3},
{8'hEE, 8'hF5, 8'hBD},
{8'hEC, 8'hF5, 8'hB8},
{8'hEE, 8'hF6, 8'hB8},
{8'hF0, 8'hF8, 8'hB9},
{8'hF1, 8'hFA, 8'hBC},
{8'hE8, 8'hF0, 8'hB8},
{8'hF3, 8'hF9, 8'hCB},
{8'hBC, 8'hC0, 8'h9D},
{8'h86, 8'h88, 8'h6F},
{8'hA8, 8'hA7, 8'hA8},
{8'h7F, 8'h7D, 8'h81},
{8'h7E, 8'h7C, 8'h7F},
{8'h7D, 8'h7B, 8'h7E},
{8'h80, 8'h7E, 8'h81},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'h7F, 8'h7D, 8'h7F},
{8'h7E, 8'h7F, 8'h77},
{8'h7E, 8'h7E, 8'h7B},
{8'h7E, 8'h7D, 8'h82},
{8'h7E, 8'h7C, 8'h88},
{8'h7E, 8'h7C, 8'h88},
{8'h7E, 8'h7D, 8'h82},
{8'h7E, 8'h7E, 8'h7C},
{8'h7C, 8'h7F, 8'h76},
{8'h86, 8'h7B, 8'h6D},
{8'hA1, 8'h64, 8'h4F},
{8'h99, 8'h6F, 8'h63},
{8'h75, 8'h7F, 8'h77},
{8'h7B, 8'h83, 8'h78},
{8'h7F, 8'h7A, 8'h88},
{8'h78, 8'h7C, 8'h94},
{8'h76, 8'h80, 8'h7B},
{8'h83, 8'h80, 8'h6A},
{8'hB5, 8'h60, 8'h52},
{8'hDA, 8'h98, 8'h73},
{8'hF6, 8'hFD, 8'hC8},
{8'hF4, 8'hF7, 8'hD3},
{8'hF9, 8'hE5, 8'hD1},
{8'hFE, 8'hFC, 8'hD7},
{8'hEB, 8'hFB, 8'hC4},
{8'hF1, 8'hED, 8'hBF},
{8'hF8, 8'hF3, 8'hC7},
{8'hF1, 8'hEB, 8'hBD},
{8'hFE, 8'hFD, 8'hCF},
{8'hFD, 8'hFC, 8'hD0},
{8'hF8, 8'hF7, 8'hCD},
{8'hFC, 8'hFC, 8'hD1},
{8'hFF, 8'hFE, 8'hD4},
{8'hFC, 8'hFC, 8'hDC},
{8'hFA, 8'hF8, 8'hD6},
{8'hE0, 8'hD1, 8'hAF},
{8'hEC, 8'hE3, 8'hBE},
{8'hF4, 8'hE6, 8'hC1},
{8'hF3, 8'hE9, 8'hC1},
{8'hF2, 8'hF1, 8'hC9},
{8'hED, 8'hEC, 8'hC4},
{8'hFC, 8'hF3, 8'hC5},
{8'hF0, 8'hE5, 8'hB7},
{8'hE5, 8'hD8, 8'hAB},
{8'hD0, 8'hBC, 8'h92},
{8'hDF, 8'hC7, 8'hA1},
{8'hB5, 8'h9E, 8'h78},
{8'hB6, 8'hB1, 8'h87},
{8'hCF, 8'hD7, 8'hAD},
{8'hA1, 8'hA7, 8'h80},
{8'h78, 8'h79, 8'h64},
{8'h79, 8'h78, 8'h73},
{8'h7A, 8'h79, 8'h74},
{8'h7B, 8'h7D, 8'h69},
{8'hCF, 8'hD3, 8'hAE},
{8'hF1, 8'hF7, 8'hCA},
{8'hEB, 8'hF1, 8'hC3},
{8'hED, 8'hF6, 8'hBA},
{8'hEF, 8'hF7, 8'hBD},
{8'hEA, 8'hF0, 8'hBC},
{8'hD2, 8'hD8, 8'hAC},
{8'hB2, 8'hB5, 8'h97},
{8'hA8, 8'hA9, 8'h9A},
{8'h9A, 8'h99, 8'h99},
{8'h7B, 8'h78, 8'h80},
{8'hFF, 8'hD7, 8'h00},
{8'h80, 8'h7E, 8'h81},
{8'h80, 8'h7E, 8'h81},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'h7F, 8'h7D, 8'h7F},
{8'h7E, 8'h7F, 8'h79},
{8'h7E, 8'h7E, 8'h7D},
{8'h7E, 8'h7D, 8'h83},
{8'h7E, 8'h7C, 8'h87},
{8'h7E, 8'h7C, 8'h87},
{8'h7E, 8'h7D, 8'h83},
{8'h7E, 8'h7E, 8'h7D},
{8'h7D, 8'h80, 8'h7B},
{8'h84, 8'h7B, 8'h74},
{8'h95, 8'h5E, 8'h4D},
{8'h91, 8'h6C, 8'h65},
{8'h78, 8'h84, 8'h82},
{8'h78, 8'h7F, 8'h76},
{8'h81, 8'h7A, 8'h87},
{8'h7E, 8'h7D, 8'h93},
{8'h82, 8'h7F, 8'h76},
{8'h87, 8'h71, 8'h57},
{8'hBC, 8'h6F, 8'h57},
{8'hF8, 8'hD0, 8'hA4},
{8'hFA, 8'hFF, 8'hCD},
{8'hEF, 8'hEE, 8'hCC},
{8'hFC, 8'hF0, 8'hD9},
{8'hFF, 8'hFE, 8'hDC},
{8'hF8, 8'hFC, 8'hCA},
{8'hF5, 8'hEE, 8'hC1},
{8'hFA, 8'hF6, 8'hCB},
{8'hE1, 8'hDC, 8'hAF},
{8'hFF, 8'hFE, 8'hD3},
{8'hFE, 8'hFD, 8'hD4},
{8'hF3, 8'hF1, 8'hC6},
{8'hEA, 8'hE7, 8'hBD},
{8'hFC, 8'hFA, 8'hD2},
{8'hFF, 8'hF6, 8'hD4},
{8'hFE, 8'hFE, 8'hD8},
{8'hF4, 8'hF1, 8'hC8},
{8'hD0, 8'hB8, 8'h90},
{8'hF8, 8'hEB, 8'hC2},
{8'hDC, 8'hD4, 8'hA7},
{8'hEE, 8'hEC, 8'hC2},
{8'hE8, 8'hD9, 8'hB3},
{8'hE0, 8'hCC, 8'h9F},
{8'hF2, 8'hE3, 8'hB4},
{8'hF7, 8'hE9, 8'hBB},
{8'hD4, 8'hBD, 8'h93},
{8'h8D, 8'h6D, 8'h46},
{8'hBC, 8'hA3, 8'h7C},
{8'hFC, 8'hF7, 8'hCB},
{8'hF5, 8'hFD, 8'hCC},
{8'hEC, 8'hF1, 8'hC4},
{8'hC6, 8'hC9, 8'hAB},
{8'hB5, 8'hB5, 8'hA9},
{8'hAA, 8'hAA, 8'h9E},
{8'hB7, 8'hBA, 8'hA0},
{8'hE3, 8'hE9, 8'hBE},
{8'hEE, 8'hF5, 8'hC3},
{8'hEF, 8'hF6, 8'hC4},
{8'hEF, 8'hF5, 8'hC6},
{8'hF1, 8'hF6, 8'hCD},
{8'hA9, 8'hAD, 8'h8C},
{8'h7E, 8'h7F, 8'h6A},
{8'h7F, 8'h80, 8'h76},
{8'h7A, 8'h79, 8'h79},
{8'h79, 8'h76, 8'h7D},
{8'h82, 8'h7F, 8'h89},
{8'h7B, 8'h79, 8'h7C},
{8'h7E, 8'h7C, 8'h7F},
{8'hFF, 8'hD7, 8'h00},
{8'h7D, 8'h7B, 8'h7E},
{8'h80, 8'h7E, 8'h81},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'h7E, 8'h7E, 8'h7D},
{8'h7E, 8'h7E, 8'h80},
{8'h7E, 8'h7D, 8'h82},
{8'h7E, 8'h7D, 8'h84},
{8'h7E, 8'h7D, 8'h84},
{8'h7D, 8'h7D, 8'h82},
{8'h7D, 8'h7D, 8'h7E},
{8'h7E, 8'h80, 8'h80},
{8'h7C, 8'h77, 8'h7A},
{8'h86, 8'h5C, 8'h52},
{8'h8D, 8'h74, 8'h72},
{8'h7A, 8'h84, 8'h87},
{8'h7D, 8'h7C, 8'h77},
{8'h86, 8'h7B, 8'h85},
{8'h83, 8'h7A, 8'h8A},
{8'h88, 8'h6F, 8'h62},
{8'hA0, 8'h6E, 8'h4D},
{8'hD5, 8'h9A, 8'h76},
{8'hFF, 8'hF6, 8'hC1},
{8'hFF, 8'hFF, 8'hCF},
{8'hEA, 8'hE0, 8'hBE},
{8'hF8, 8'hF7, 8'hDB},
{8'hFB, 8'hFF, 8'hDC},
{8'hFF, 8'hF9, 8'hD2},
{8'hF9, 8'hF5, 8'hCC},
{8'hFD, 8'hF8, 8'hCF},
{8'hD6, 8'hD1, 8'hA8},
{8'hF2, 8'hEE, 8'hC6},
{8'hFF, 8'hFC, 8'hD3},
{8'hFE, 8'hFC, 8'hD3},
{8'hE2, 8'hDD, 8'hB3},
{8'hE2, 8'hDC, 8'hB4},
{8'hFF, 8'hF6, 8'hD4},
{8'hFB, 8'hFA, 8'hD0},
{8'hFD, 8'hFF, 8'hCF},
{8'hEB, 8'hD3, 8'hA3},
{8'hCD, 8'hB1, 8'h81},
{8'hEF, 8'hE9, 8'hB5},
{8'hBE, 8'hAE, 8'h7E},
{8'hF4, 8'hD5, 8'hB2},
{8'hE0, 8'hC8, 8'h9B},
{8'hE8, 8'hD5, 8'hA6},
{8'hF2, 8'hE1, 8'hB2},
{8'hF3, 8'hDA, 8'hAE},
{8'h92, 8'h70, 8'h49},
{8'hAF, 8'h94, 8'h6E},
{8'hDD, 8'hD1, 8'hA5},
{8'hF1, 8'hF4, 8'hC2},
{8'hF0, 8'hF7, 8'hC1},
{8'hF0, 8'hF3, 8'hCE},
{8'hEC, 8'hED, 8'hDA},
{8'hF5, 8'hF6, 8'hE4},
{8'hD5, 8'hD9, 8'hB8},
{8'hD3, 8'hD9, 8'hA9},
{8'hF4, 8'hFB, 8'hC5},
{8'hEF, 8'hF7, 8'hC2},
{8'hF5, 8'hF9, 8'hD6},
{8'hC5, 8'hC7, 8'hAE},
{8'h7A, 8'h7A, 8'h6E},
{8'h7D, 8'h7B, 8'h7C},
{8'h84, 8'h82, 8'h8A},
{8'h80, 8'h7D, 8'h86},
{8'h7F, 8'h7D, 8'h82},
{8'h7C, 8'h7A, 8'h7D},
{8'h81, 8'h7F, 8'h81},
{8'h7F, 8'h7D, 8'h7F},
{8'h80, 8'h7E, 8'h81},
{8'h83, 8'h81, 8'h84},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'h7E, 8'h7D, 8'h81},
{8'h7D, 8'h7D, 8'h7F},
{8'h7D, 8'h7D, 8'h7E},
{8'h7D, 8'h7D, 8'h7C},
{8'h7E, 8'h7E, 8'h7E},
{8'h80, 8'h80, 8'h81},
{8'h85, 8'h84, 8'h86},
{8'h7B, 8'h7C, 8'h82},
{8'h72, 8'h71, 8'h7B},
{8'h7C, 8'h60, 8'h58},
{8'h8B, 8'h7E, 8'h7F},
{8'h78, 8'h7F, 8'h89},
{8'h84, 8'h7D, 8'h7B},
{8'h8A, 8'h7E, 8'h83},
{8'h85, 8'h75, 8'h7C},
{8'h90, 8'h61, 8'h4D},
{8'hBD, 8'h74, 8'h4A},
{8'hEA, 8'hC4, 8'h93},
{8'hFD, 8'hFF, 8'hC6},
{8'hFD, 8'hFD, 8'hCE},
{8'hE6, 8'hD2, 8'hB0},
{8'hF7, 8'hF7, 8'hD7},
{8'hF2, 8'hFE, 8'hD9},
{8'hFF, 8'hEE, 8'hD3},
{8'hFD, 8'hFA, 8'hD2},
{8'hFD, 8'hFD, 8'hD7},
{8'hE6, 8'hE1, 8'hBA},
{8'hCF, 8'hC5, 8'h9C},
{8'hFD, 8'hF7, 8'hCE},
{8'hFE, 8'hF9, 8'hD0},
{8'hFB, 8'hF7, 8'hCD},
{8'hC1, 8'hB4, 8'h89},
{8'hF1, 8'hD7, 8'hB2},
{8'hF4, 8'hF4, 8'hC0},
{8'hF9, 8'hFD, 8'hC4},
{8'hF9, 8'hE5, 8'hB0},
{8'hC1, 8'hA2, 8'h6D},
{8'hD9, 8'hD0, 8'h96},
{8'hD7, 8'hC0, 8'h8E},
{8'hC6, 8'h86, 8'h65},
{8'hF6, 8'hD8, 8'hAC},
{8'hF9, 8'hE7, 8'hB7},
{8'hFD, 8'hF2, 8'hC1},
{8'hFD, 8'hEC, 8'hBE},
{8'hCA, 8'hA7, 8'h7D},
{8'hC6, 8'hAC, 8'h84},
{8'hD8, 8'hC7, 8'h9B},
{8'hE0, 8'hDC, 8'hAB},
{8'hF1, 8'hF9, 8'hBD},
{8'hED, 8'hF3, 8'hC6},
{8'hEA, 8'hEB, 8'hD2},
{8'hD4, 8'hD6, 8'hC0},
{8'hB9, 8'hBD, 8'h9A},
{8'hDE, 8'hE5, 8'hB2},
{8'hED, 8'hF5, 8'hBC},
{8'hEF, 8'hF6, 8'hC0},
{8'hDF, 8'hE3, 8'hC1},
{8'h81, 8'h83, 8'h6E},
{8'h7B, 8'h7A, 8'h73},
{8'h7E, 8'h7B, 8'h81},
{8'h7B, 8'h78, 8'h81},
{8'h80, 8'h7D, 8'h81},
{8'h8C, 8'h8B, 8'h84},
{8'h79, 8'h7A, 8'h6D},
{8'h85, 8'h83, 8'h85},
{8'h91, 8'h8F, 8'h92},
{8'h8D, 8'h8B, 8'h8E},
{8'h80, 8'h7E, 8'h81},
{8'h7E, 8'h7C, 8'h7F},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'h80, 8'h7E, 8'h81},
{8'h7F, 8'h7E, 8'h83},
{8'h7C, 8'h7C, 8'h7E},
{8'h86, 8'h87, 8'h80},
{8'h7F, 8'h81, 8'h76},
{8'h7B, 8'h7D, 8'h71},
{8'hB0, 8'hB2, 8'hAB},
{8'hE6, 8'hE5, 8'hE6},
{8'h94, 8'h94, 8'h9B},
{8'h71, 8'h6F, 8'h7A},
{8'h78, 8'h68, 8'h5F},
{8'h82, 8'h81, 8'h82},
{8'h77, 8'h7B, 8'h87},
{8'h85, 8'h76, 8'h75},
{8'h82, 8'h78, 8'h76},
{8'h7C, 8'h68, 8'h67},
{8'hA1, 8'h60, 8'h45},
{8'hCE, 8'h7D, 8'h49},
{8'hF7, 8'hD6, 8'h9E},
{8'hF9, 8'hFF, 8'hCB},
{8'hF7, 8'hF6, 8'hC8},
{8'hD3, 8'hB3, 8'h93},
{8'hF6, 8'hF7, 8'hD0},
{8'hF5, 8'hFE, 8'hD8},
{8'hFD, 8'hE3, 8'hCA},
{8'hFC, 8'hF8, 8'hD1},
{8'hFF, 8'hFF, 8'hD6},
{8'hFA, 8'hF6, 8'hCD},
{8'hB0, 8'h9D, 8'h75},
{8'hE7, 8'hDA, 8'hB1},
{8'hEC, 8'hDC, 8'hB2},
{8'hFF, 8'hFC, 8'hD1},
{8'hE6, 8'hD7, 8'hA9},
{8'hBD, 8'h93, 8'h6C},
{8'hE9, 8'hDD, 8'hAA},
{8'hE7, 8'hE0, 8'hA5},
{8'hFF, 8'hF5, 8'hBC},
{8'hD2, 8'hB2, 8'h7A},
{8'hB0, 8'h97, 8'h5E},
{8'hF6, 8'hDF, 8'hAE},
{8'hB1, 8'h6D, 8'h48},
{8'hB4, 8'h8A, 8'h5E},
{8'hE4, 8'hC8, 8'h98},
{8'hFC, 8'hEB, 8'hBA},
{8'hFC, 8'hEE, 8'hBE},
{8'hF4, 8'hE3, 8'hB8},
{8'hA8, 8'h85, 8'h5B},
{8'hA4, 8'h8A, 8'h5D},
{8'hEF, 8'hE7, 8'hB5},
{8'hF3, 8'hF8, 8'hBD},
{8'hED, 8'hF4, 8'hC7},
{8'hF3, 8'hF4, 8'hDC},
{8'hC8, 8'hCA, 8'hB4},
{8'hD1, 8'hD5, 8'hB3},
{8'hED, 8'hF3, 8'hC3},
{8'hE9, 8'hF0, 8'hBC},
{8'hF2, 8'hF9, 8'hC7},
{8'hD3, 8'hD7, 8'hB4},
{8'h9B, 8'h9E, 8'h82},
{8'h94, 8'h95, 8'h85},
{8'h89, 8'h88, 8'h80},
{8'h8C, 8'h8B, 8'h85},
{8'hA4, 8'hA5, 8'h98},
{8'hA4, 8'hA5, 8'h91},
{8'hA7, 8'hAA, 8'h92},
{8'hA0, 8'h9E, 8'h9F},
{8'h8B, 8'h89, 8'h8C},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'h7B, 8'h7B, 8'h7F},
{8'h9B, 8'h9B, 8'h98},
{8'hE3, 8'hE5, 8'hD5},
{8'hB7, 8'hBB, 8'hA3},
{8'h76, 8'h7A, 8'h62},
{8'hBB, 8'hBE, 8'hAE},
{8'hFF, 8'hFF, 8'hFC},
{8'hDB, 8'hDB, 8'hE0},
{8'h86, 8'h81, 8'h88},
{8'h76, 8'h6E, 8'h5E},
{8'h73, 8'h7A, 8'h74},
{8'h76, 8'h78, 8'h82},
{8'h99, 8'h86, 8'h82},
{8'hAA, 8'hA4, 8'h9C},
{8'h8C, 8'h7A, 8'h70},
{8'hAD, 8'h61, 8'h40},
{8'hCF, 8'h87, 8'h48},
{8'hEF, 8'hD3, 8'h99},
{8'hF9, 8'hFD, 8'hCF},
{8'hF6, 8'hF7, 8'hCE},
{8'hC2, 8'h9A, 8'h78},
{8'hF7, 8'hEF, 8'hC0},
{8'hFB, 8'hFF, 8'hD5},
{8'hF1, 8'hDD, 8'hBF},
{8'hF6, 8'hF3, 8'hC9},
{8'hFE, 8'hFA, 8'hCF},
{8'hFF, 8'hFE, 8'hD4},
{8'hCD, 8'hB8, 8'h8E},
{8'hC6, 8'hA6, 8'h7C},
{8'hEB, 8'hD5, 8'hA8},
{8'hE5, 8'hCC, 8'h9C},
{8'hFF, 8'hF6, 8'hC4},
{8'hCA, 8'hAA, 8'h7E},
{8'hBE, 8'h97, 8'h6B},
{8'hDD, 8'hBB, 8'h89},
{8'hF1, 8'hDD, 8'hA5},
{8'hDF, 8'hC0, 8'h88},
{8'hA6, 8'h73, 8'h41},
{8'hDC, 8'hB0, 8'h83},
{8'hDF, 8'hAD, 8'h82},
{8'hA0, 8'h6E, 8'h40},
{8'hA6, 8'h7F, 8'h4D},
{8'hD3, 8'hBB, 8'h88},
{8'hE9, 8'hD0, 8'h9F},
{8'hF5, 8'hDE, 8'hB1},
{8'hBF, 8'hA0, 8'h75},
{8'h96, 8'h75, 8'h47},
{8'hFA, 8'hEA, 8'hB8},
{8'hEC, 8'hF2, 8'hBA},
{8'hED, 8'hF3, 8'hCB},
{8'hF5, 8'hF6, 8'hE3},
{8'hF1, 8'hF1, 8'hE3},
{8'hF1, 8'hF3, 8'hD9},
{8'hED, 8'hF2, 8'hCB},
{8'hEF, 8'hF5, 8'hC9},
{8'hE6, 8'hEB, 8'hC2},
{8'hA5, 8'hA8, 8'h89},
{8'h9E, 8'hA1, 8'h84},
{8'hA7, 8'hAA, 8'h8E},
{8'hB3, 8'hB6, 8'h9B},
{8'hC9, 8'hCB, 8'hB3},
{8'hAD, 8'hAF, 8'h98},
{8'hE8, 8'hEA, 8'hD3},
{8'hAA, 8'hAC, 8'h98},
{8'h79, 8'h77, 8'h78},
{8'h7D, 8'h7B, 8'h7F},
{8'h7C, 8'h7A, 8'h7D},
{8'h80, 8'h7E, 8'h81},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'h80, 8'h7E, 8'h80},
{8'h7D, 8'h7C, 8'h7D},
{8'h9A, 8'h9B, 8'h92},
{8'hED, 8'hF0, 8'hD7},
{8'hEC, 8'hF2, 8'hCF},
{8'hAD, 8'hB3, 8'h8F},
{8'hB6, 8'hB9, 8'hA2},
{8'hFC, 8'hFD, 8'hF4},
{8'hFE, 8'hFD, 8'hFE},
{8'hC6, 8'hBD, 8'hBE},
{8'h9D, 8'h99, 8'h7F},
{8'hAA, 8'hB7, 8'hAA},
{8'hB6, 8'hB6, 8'hBD},
{8'hEE, 8'hE0, 8'hDA},
{8'hD3, 8'hD1, 8'hC3},
{8'hCA, 8'hBA, 8'hA9},
{8'hB8, 8'h66, 8'h3E},
{8'hCA, 8'h91, 8'h4A},
{8'hDE, 8'hC6, 8'h8F},
{8'hF7, 8'hF6, 8'hD0},
{8'hF7, 8'hF7, 8'hD4},
{8'hC5, 8'h94, 8'h71},
{8'hF6, 8'hDC, 8'hAB},
{8'hFF, 8'hFF, 8'hD4},
{8'hEB, 8'hE7, 8'hC0},
{8'hE3, 8'hE3, 8'hB4},
{8'hFC, 8'hF5, 8'hC8},
{8'hF4, 8'hE8, 8'hBB},
{8'hED, 8'hD4, 8'hA8},
{8'hBF, 8'h92, 8'h64},
{8'hE6, 8'hC1, 8'h90},
{8'hC8, 8'hA3, 8'h6E},
{8'hE4, 8'hC8, 8'h90},
{8'hEC, 8'hD8, 8'hA8},
{8'hCE, 8'h8E, 8'h6B},
{8'hD9, 8'h96, 8'h6F},
{8'hCD, 8'hB0, 8'h79},
{8'hEC, 8'hD3, 8'h9C},
{8'hB4, 8'h6A, 8'h41},
{8'hB4, 8'h70, 8'h48},
{8'hED, 8'hD8, 8'hA6},
{8'hC5, 8'h94, 8'h66},
{8'hA9, 8'h7C, 8'h4A},
{8'hA0, 8'h7E, 8'h4A},
{8'hB0, 8'h8E, 8'h5C},
{8'hCE, 8'hA4, 8'h76},
{8'hC7, 8'h9B, 8'h6F},
{8'h89, 8'h65, 8'h37},
{8'hE8, 8'hD3, 8'hA2},
{8'hF2, 8'hF8, 8'hC5},
{8'hE7, 8'hEB, 8'hCA},
{8'hF2, 8'hF3, 8'hE7},
{8'hF7, 8'hF7, 8'hF1},
{8'hEA, 8'hEB, 8'hDB},
{8'hE2, 8'hE5, 8'hC9},
{8'hE7, 8'hEB, 8'hCA},
{8'hDD, 8'hE1, 8'hC3},
{8'hA2, 8'hA3, 8'h93},
{8'h7E, 8'h7F, 8'h6A},
{8'hA2, 8'hA6, 8'h88},
{8'hBA, 8'hBE, 8'h9A},
{8'h95, 8'h99, 8'h78},
{8'hD4, 8'hD5, 8'hC0},
{8'hF9, 8'hF9, 8'hEF},
{8'hAF, 8'hAE, 8'hAD},
{8'h75, 8'h73, 8'h76},
{8'h7E, 8'h7C, 8'h7F},
{8'h80, 8'h7E, 8'h81},
{8'h7D, 8'h7B, 8'h7E},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'h7F, 8'h7D, 8'h7F},
{8'h7F, 8'h7D, 8'h7F},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'h7F, 8'h7D, 8'h81},
{8'h7F, 8'h7D, 8'h82},
{8'h7F, 8'h7C, 8'h83},
{8'h7E, 8'h7C, 8'h83},
{8'h7B, 8'h7B, 8'h7A},
{8'h82, 8'h85, 8'h77},
{8'hDA, 8'hDF, 8'hC1},
{8'hED, 8'hF5, 8'hC9},
{8'hDE, 8'hE6, 8'hBB},
{8'hD5, 8'hD9, 8'hBC},
{8'hF9, 8'hFA, 8'hF0},
{8'hFA, 8'hF9, 8'hFA},
{8'hF4, 8'hE9, 8'hE7},
{8'hD4, 8'hD3, 8'hBA},
{8'hEA, 8'hF8, 8'hEA},
{8'hF7, 8'hF6, 8'hFA},
{8'hFF, 8'hF6, 8'hEE},
{8'hBE, 8'hC0, 8'hB0},
{8'h96, 8'h86, 8'h74},
{8'hAC, 8'h5A, 8'h32},
{8'hCC, 8'h96, 8'h4F},
{8'hD7, 8'hB7, 8'h82},
{8'hF4, 8'hEE, 8'hC6},
{8'hF7, 8'hF6, 8'hD1},
{8'hCD, 8'h97, 8'h74},
{8'hE7, 8'hC2, 8'h93},
{8'hFD, 8'hFD, 8'hC9},
{8'hE9, 8'hF3, 8'hC2},
{8'hCD, 8'hC8, 8'h96},
{8'hFE, 8'hFA, 8'hC9},
{8'hDA, 8'hBF, 8'h8F},
{8'hF7, 8'hE1, 8'hB3},
{8'hCA, 8'h9D, 8'h6B},
{8'hBC, 8'h8B, 8'h56},
{8'hD8, 8'hA9, 8'h71},
{8'hB5, 8'h92, 8'h55},
{8'hE1, 8'hD4, 8'h9F},
{8'hFC, 8'hB6, 8'h95},
{8'hE5, 8'h90, 8'h72},
{8'hB2, 8'h89, 8'h58},
{8'hD9, 8'hB9, 8'h86},
{8'hC7, 8'h73, 8'h4F},
{8'h9C, 8'h51, 8'h2A},
{8'hD5, 8'hC6, 8'h8E},
{8'hED, 8'hCE, 8'h9D},
{8'hBB, 8'h8C, 8'h5B},
{8'hE7, 8'hCC, 8'h97},
{8'hE9, 8'hD6, 8'hA3},
{8'hDE, 8'hC2, 8'h93},
{8'hC9, 8'h9F, 8'h73},
{8'hA2, 8'h7B, 8'h4D},
{8'hD9, 8'hC1, 8'h90},
{8'hED, 8'hF0, 8'hC3},
{8'hE7, 8'hEA, 8'hCF},
{8'hF2, 8'hF1, 8'hEA},
{8'hFB, 8'hFA, 8'hF8},
{8'hF0, 8'hF0, 8'hE6},
{8'hE1, 8'hE2, 8'hCE},
{8'hE2, 8'hE4, 8'hCC},
{8'hEB, 8'hED, 8'hD7},
{8'hEE, 8'hEC, 8'hE8},
{8'hDD, 8'hDD, 8'hD1},
{8'hEB, 8'hED, 8'hD3},
{8'hDE, 8'hE1, 8'hBE},
{8'hD7, 8'hDB, 8'hB9},
{8'hF8, 8'hF8, 8'hE6},
{8'hFA, 8'hF9, 8'hF5},
{8'hC6, 8'hC2, 8'hC8},
{8'h7E, 8'h7D, 8'h7D},
{8'h7F, 8'h7D, 8'h7C},
{8'h7D, 8'h7B, 8'h7D},
{8'h82, 8'h80, 8'h83},
{8'h81, 8'h7F, 8'h82},
{8'h7F, 8'h7D, 8'h81},
{8'h7E, 8'h7C, 8'h7F},
{8'h7F, 8'h7D, 8'h7F},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'h7E, 8'h7E, 8'h7E},
{8'h7E, 8'h7E, 8'h7D},
{8'h7E, 8'h7E, 8'h7E},
{8'h7E, 8'h7E, 8'h7F},
{8'h7B, 8'h7A, 8'h80},
{8'h7E, 8'h7C, 8'h87},
{8'h7D, 8'h7A, 8'h8B},
{8'h78, 8'h76, 8'h87},
{8'h77, 8'h7C, 8'h7C},
{8'h78, 8'h80, 8'h6F},
{8'hC6, 8'hD0, 8'hAA},
{8'hEA, 8'hF5, 8'hC0},
{8'hE4, 8'hEE, 8'hBC},
{8'hEC, 8'hF1, 8'hD2},
{8'hFA, 8'hFA, 8'hF4},
{8'hF8, 8'hF3, 8'hFB},
{8'hF9, 8'hEE, 8'hE9},
{8'hDF, 8'hDF, 8'hEA},
{8'hED, 8'hF0, 8'hFC},
{8'hF8, 8'hF1, 8'hEF},
{8'hFE, 8'hFB, 8'hF1},
{8'h9F, 8'h9E, 8'h9A},
{8'h81, 8'h63, 8'h59},
{8'hA9, 8'h5D, 8'h41},
{8'hE1, 8'h8C, 8'h5E},
{8'hD0, 8'hA7, 8'h6D},
{8'hE2, 8'hDD, 8'h9F},
{8'hF9, 8'hF1, 8'hBA},
{8'hD5, 8'hA3, 8'h7C},
{8'hD6, 8'h9E, 8'h7D},
{8'hF6, 8'hE5, 8'hB9},
{8'hF4, 8'hF9, 8'hC4},
{8'hD4, 8'hAE, 8'h7D},
{8'hF4, 8'hEA, 8'hB3},
{8'hDF, 8'hBB, 8'h87},
{8'hDD, 8'hA7, 8'h72},
{8'hCD, 8'hA7, 8'h69},
{8'hEA, 8'hB5, 8'h78},
{8'hE4, 8'h9D, 8'h67},
{8'hBF, 8'h8C, 8'h4D},
{8'hB0, 8'h82, 8'h40},
{8'hE1, 8'hAB, 8'h7C},
{8'hF4, 8'hB7, 8'h9F},
{8'hBD, 8'h70, 8'h5E},
{8'hC4, 8'h77, 8'h5A},
{8'hC7, 8'h7D, 8'h53},
{8'h8C, 8'h47, 8'h17},
{8'hC7, 8'h8E, 8'h5C},
{8'hFF, 8'hF7, 8'hBC},
{8'hC7, 8'hA7, 8'h74},
{8'hDC, 8'hBD, 8'h8D},
{8'hF2, 8'hE3, 8'hB0},
{8'hF9, 8'hED, 8'hBD},
{8'hEE, 8'hCD, 8'hA7},
{8'h9B, 8'h70, 8'h43},
{8'hBF, 8'hB8, 8'h7F},
{8'hEB, 8'hEC, 8'hC6},
{8'hEF, 8'hEE, 8'hD2},
{8'hF5, 8'hF1, 8'hE2},
{8'hFE, 8'hFB, 8'hF5},
{8'hFA, 8'hF5, 8'hF2},
{8'hE3, 8'hDF, 8'hD6},
{8'hE1, 8'hDE, 8'hCD},
{8'hEB, 8'hE9, 8'hD4},
{8'hF0, 8'hE9, 8'hE6},
{8'hFB, 8'hF6, 8'hF0},
{8'hF8, 8'hF6, 8'hE8},
{8'hF0, 8'hF1, 8'hDC},
{8'hED, 8'hEF, 8'hD5},
{8'hF4, 8'hF4, 8'hDB},
{8'hFB, 8'hF9, 8'hE1},
{8'hF6, 8'hF2, 8'hDC},
{8'hB2, 8'hB5, 8'h97},
{8'h7A, 8'h7B, 8'h66},
{8'h80, 8'h7F, 8'h77},
{8'h84, 8'h82, 8'h85},
{8'h7D, 8'h7A, 8'h83},
{8'h7F, 8'h7C, 8'h84},
{8'h7F, 8'h7D, 8'h7E},
{8'h7E, 8'h7D, 8'h79},
{8'h80, 8'h7E, 8'h80},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'h7E, 8'h7C, 8'h85},
{8'h7E, 8'h7D, 8'h83},
{8'h7E, 8'h7E, 8'h7F},
{8'h7E, 8'h7F, 8'h79},
{8'h82, 8'h84, 8'h79},
{8'h8A, 8'h8D, 8'h7E},
{8'h85, 8'h88, 8'h76},
{8'h8D, 8'h90, 8'h7E},
{8'h8B, 8'h8E, 8'h8B},
{8'h7B, 8'h80, 8'h74},
{8'hB1, 8'hB6, 8'h9B},
{8'hE7, 8'hEC, 8'hC7},
{8'hE4, 8'hE8, 8'hC3},
{8'hEF, 8'hF0, 8'hD6},
{8'hFA, 8'hF9, 8'hEC},
{8'hFA, 8'hF6, 8'hF0},
{8'hFC, 8'hF4, 8'hD5},
{8'hE5, 8'hE6, 8'hDD},
{8'hEB, 8'hED, 8'hF2},
{8'hFE, 8'hF3, 8'hF0},
{8'hDA, 8'hD4, 8'hCB},
{8'h6E, 8'h6C, 8'h69},
{8'h89, 8'h6C, 8'h60},
{8'hAB, 8'h62, 8'h41},
{8'hD7, 8'h85, 8'h56},
{8'hC7, 8'h93, 8'h5B},
{8'hCE, 8'hB8, 8'h7B},
{8'hFE, 8'hF3, 8'hBA},
{8'hE2, 8'hB4, 8'h86},
{8'hD6, 8'h9E, 8'h75},
{8'hE3, 8'hBD, 8'h90},
{8'hF7, 8'hE9, 8'hB6},
{8'hCF, 8'hBE, 8'h8B},
{8'hCC, 8'hB0, 8'h7F},
{8'hF6, 8'hE0, 8'hAC},
{8'hB1, 8'h86, 8'h51},
{8'hDB, 8'hA4, 8'h75},
{8'hF5, 8'hC0, 8'h92},
{8'hF9, 8'hC0, 8'h93},
{8'hC8, 8'h82, 8'h5A},
{8'h9D, 8'h59, 8'h2E},
{8'h8B, 8'h53, 8'h34},
{8'h92, 8'h62, 8'h51},
{8'h91, 8'h59, 8'h4C},
{8'h82, 8'h3D, 8'h27},
{8'hB1, 8'h67, 8'h42},
{8'h93, 8'h4F, 8'h23},
{8'hAD, 8'h78, 8'h48},
{8'hFF, 8'hF9, 8'hC3},
{8'hE7, 8'hCF, 8'h9E},
{8'hCB, 8'hAB, 8'h7C},
{8'hC6, 8'hB3, 8'h80},
{8'hC8, 8'hA7, 8'h78},
{8'hAF, 8'h73, 8'h4D},
{8'h81, 8'h53, 8'h26},
{8'hD8, 8'hCE, 8'h97},
{8'hF3, 8'hF3, 8'hD0},
{8'hED, 8'hEC, 8'hD3},
{8'hFE, 8'hFC, 8'hED},
{8'hFD, 8'hF8, 8'hF2},
{8'hFE, 8'hFA, 8'hF5},
{8'hEF, 8'hEB, 8'hE2},
{8'hE3, 8'hE0, 8'hCF},
{8'hF3, 8'hF1, 8'hDC},
{8'hF7, 8'hF3, 8'hEC},
{8'hFC, 8'hF9, 8'hF3},
{8'hFC, 8'hFB, 8'hF3},
{8'hF5, 8'hF5, 8'hEA},
{8'hF0, 8'hF0, 8'hE2},
{8'hF6, 8'hF6, 8'hE6},
{8'hF9, 8'hF7, 8'hE7},
{8'hF3, 8'hF2, 8'hDF},
{8'hE7, 8'hE9, 8'hCE},
{8'h9E, 8'hA0, 8'h8C},
{8'h7A, 8'h7A, 8'h72},
{8'h78, 8'h76, 8'h79},
{8'h7E, 8'h7B, 8'h84},
{8'h7D, 8'h7A, 8'h81},
{8'h7E, 8'h7C, 8'h7D},
{8'h7E, 8'h7D, 8'h79},
{8'h7F, 8'h7D, 8'h7F},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'h7F, 8'h7D, 8'h81},
{8'h7E, 8'h7C, 8'h89},
{8'h7E, 8'h7C, 8'h87},
{8'h7E, 8'h7E, 8'h80},
{8'h7A, 8'h7B, 8'h72},
{8'h94, 8'h97, 8'h80},
{8'hE0, 8'hE6, 8'hC2},
{8'hE8, 8'hEF, 8'hC1},
{8'hEA, 8'hF1, 8'hC1},
{8'hE2, 8'hE1, 8'hDA},
{8'hE3, 8'hE3, 8'hDD},
{8'hEE, 8'hEC, 8'hE2},
{8'hFA, 8'hF8, 8'hE9},
{8'hF4, 8'hF2, 8'hE0},
{8'hF1, 8'hED, 8'hD9},
{8'hEF, 8'hEC, 8'hD6},
{8'hFC, 8'hF8, 8'hDC},
{8'hF6, 8'hEC, 8'hA8},
{8'hEB, 8'hEC, 8'hC7},
{8'hED, 8'hED, 8'hE2},
{8'hFE, 8'hEF, 8'hE6},
{8'hD2, 8'hC7, 8'hC1},
{8'h93, 8'h90, 8'h8F},
{8'h92, 8'h77, 8'h69},
{8'hA4, 8'h60, 8'h3A},
{8'hC1, 8'h75, 8'h45},
{8'hBF, 8'h7C, 8'h4A},
{8'hBE, 8'h8A, 8'h54},
{8'hFC, 8'hEB, 8'hB1},
{8'hDE, 8'hB8, 8'h7F},
{8'hCF, 8'h9D, 8'h6A},
{8'hC1, 8'h83, 8'h55},
{8'hD3, 8'h9B, 8'h6F},
{8'hEC, 8'hDC, 8'hA6},
{8'hAB, 8'h7A, 8'h4B},
{8'hEF, 8'hD6, 8'hA2},
{8'hC4, 8'hA3, 8'h6E},
{8'hCB, 8'h7D, 8'h59},
{8'hE5, 8'hA8, 8'h87},
{8'hF4, 8'hCD, 8'hAB},
{8'hBF, 8'h71, 8'h5E},
{8'hA2, 8'h5B, 8'h48},
{8'h60, 8'h3F, 8'h2F},
{8'h38, 8'h37, 8'h28},
{8'h91, 8'h86, 8'h78},
{8'hBF, 8'h90, 8'h7E},
{8'h8E, 8'h41, 8'h27},
{8'h9C, 8'h54, 8'h2F},
{8'hBC, 8'h8A, 8'h5D},
{8'hFE, 8'hFC, 8'hCC},
{8'hF8, 8'hEA, 8'hBD},
{8'hDC, 8'hC1, 8'h94},
{8'hE1, 8'hCE, 8'h9D},
{8'hAF, 8'h8A, 8'h5E},
{8'h88, 8'h49, 8'h25},
{8'h99, 8'h66, 8'h3E},
{8'hF7, 8'hED, 8'hB9},
{8'hF0, 8'hEE, 8'hD1},
{8'hE5, 8'hE2, 8'hCD},
{8'hF6, 8'hF2, 8'hE4},
{8'hFE, 8'hFA, 8'hF2},
{8'hFB, 8'hF7, 8'hF0},
{8'hFD, 8'hF9, 8'hEF},
{8'hF3, 8'hF0, 8'hDF},
{8'hEF, 8'hEE, 8'hD9},
{8'hF8, 8'hF9, 8'hEC},
{8'hFA, 8'hFA, 8'hF2},
{8'hFB, 8'hFA, 8'hF5},
{8'hF9, 8'hF8, 8'hF6},
{8'hF5, 8'hF3, 8'hF2},
{8'hF8, 8'hF7, 8'hF3},
{8'hF7, 8'hF8, 8'hF0},
{8'hEE, 8'hF0, 8'hE3},
{8'hCC, 8'hCE, 8'hB8},
{8'h80, 8'h82, 8'h71},
{8'h93, 8'h92, 8'h8C},
{8'hB5, 8'hB3, 8'hB6},
{8'hD8, 8'hD5, 8'hDC},
{8'h9D, 8'h9B, 8'hA1},
{8'h7C, 8'h7A, 8'h7C},
{8'h7E, 8'h7D, 8'h7B},
{8'h7F, 8'h7D, 8'h7F},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'h7E, 8'h7D, 8'h85},
{8'h7E, 8'h7D, 8'h84},
{8'h7E, 8'h7E, 8'h80},
{8'h7D, 8'h7E, 8'h79},
{8'h81, 8'h83, 8'h73},
{8'hB1, 8'hB5, 8'h99},
{8'hC7, 8'hCE, 8'hA6},
{8'hD5, 8'hDB, 8'hB1},
{8'hF5, 8'hF3, 8'hE6},
{8'hFE, 8'hFB, 8'hF5},
{8'hFD, 8'hF9, 8'hF8},
{8'hFA, 8'hF3, 8'hF5},
{8'hFB, 8'hF4, 8'hF0},
{8'hFB, 8'hF5, 8'hE5},
{8'hEF, 8'hEA, 8'hCE},
{8'hEF, 8'hEA, 8'hBF},
{8'hE1, 8'hD8, 8'h7C},
{8'hEA, 8'hED, 8'hB4},
{8'hF1, 8'hEF, 8'hD9},
{8'hF8, 8'hE6, 8'hD9},
{8'hFD, 8'hF2, 8'hEB},
{8'hE2, 8'hE3, 8'hE2},
{8'hDF, 8'hCB, 8'hBC},
{8'h9C, 8'h60, 8'h39},
{8'hB1, 8'h6A, 8'h3C},
{8'hB7, 8'h69, 8'h3C},
{8'hAE, 8'h5E, 8'h2F},
{8'hF2, 8'hC2, 8'h8B},
{8'hD7, 8'hB3, 8'h76},
{8'hDD, 8'hB3, 8'h79},
{8'hC9, 8'h80, 8'h55},
{8'hD6, 8'h76, 8'h55},
{8'hEE, 8'hC3, 8'h8F},
{8'hB5, 8'h76, 8'h44},
{8'hCF, 8'h95, 8'h60},
{8'hE2, 8'hB2, 8'h7D},
{8'hE3, 8'h97, 8'h6D},
{8'hCA, 8'h8A, 8'h67},
{8'hCF, 8'hA5, 8'h87},
{8'hDA, 8'hA5, 8'h93},
{8'h9E, 8'h80, 8'h75},
{8'h16, 8'h20, 8'h11},
{8'h0C, 8'h34, 8'h22},
{8'h29, 8'h4C, 8'h3B},
{8'hDC, 8'hC8, 8'hB7},
{8'h85, 8'h3B, 8'h26},
{8'h9F, 8'h4E, 8'h2F},
{8'hC5, 8'h8C, 8'h65},
{8'hF7, 8'hF8, 8'hCA},
{8'hFE, 8'hF6, 8'hCC},
{8'hE9, 8'hD4, 8'hAA},
{8'hE6, 8'hD7, 8'hA7},
{8'hBF, 8'h99, 8'h6E},
{8'h94, 8'h51, 8'h31},
{8'hAF, 8'h7C, 8'h59},
{8'hDF, 8'hD1, 8'hA5},
{8'hF2, 8'hF0, 8'hD9},
{8'hF4, 8'hF2, 8'hE0},
{8'hFB, 8'hF7, 8'hEB},
{8'hFF, 8'hFC, 8'hF3},
{8'hFE, 8'hFC, 8'hF4},
{8'hFC, 8'hF9, 8'hED},
{8'hFB, 8'hF9, 8'hE9},
{8'hF4, 8'hF2, 8'hDE},
{8'hF3, 8'hF6, 8'hE7},
{8'hF5, 8'hF7, 8'hEC},
{8'hF9, 8'hF7, 8'hF1},
{8'hFB, 8'hF6, 8'hF5},
{8'hFA, 8'hF6, 8'hF5},
{8'hFC, 8'hF9, 8'hF8},
{8'hF7, 8'hF8, 8'hF3},
{8'hEC, 8'hEE, 8'hE7},
{8'hEF, 8'hEF, 8'hE0},
{8'hE8, 8'hE7, 8'hDC},
{8'hEF, 8'hEE, 8'hEA},
{8'hF5, 8'hF3, 8'hF5},
{8'hF9, 8'hF6, 8'hFB},
{8'hA3, 8'hA1, 8'hA6},
{8'h7D, 8'h7B, 8'h7D},
{8'h80, 8'h7E, 8'h7F},
{8'h7F, 8'h7D, 8'h7F},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'h7F, 8'h80, 8'h7C},
{8'h7F, 8'h80, 8'h7F},
{8'h80, 8'h80, 8'h83},
{8'h82, 8'h81, 8'h86},
{8'h83, 8'h83, 8'h85},
{8'h78, 8'h79, 8'h75},
{8'h7C, 8'h7E, 8'h74},
{8'h9F, 8'hA1, 8'h90},
{8'hD5, 8'hD5, 8'hBC},
{8'hF5, 8'hF3, 8'hE3},
{8'hFC, 8'hF9, 8'hF5},
{8'hFB, 8'hF4, 8'hF7},
{8'hF8, 8'hF1, 8'hF1},
{8'hFF, 8'hF8, 8'hEB},
{8'hF9, 8'hF4, 8'hD9},
{8'hEA, 8'hE5, 8'hBA},
{8'hE0, 8'hD6, 8'h7B},
{8'hE9, 8'hEB, 8'hB2},
{8'hF7, 8'hF4, 8'hDC},
{8'hFC, 8'hEC, 8'hDB},
{8'hFD, 8'hF4, 8'hEA},
{8'hE7, 8'hEA, 8'hEA},
{8'hD9, 8'hCC, 8'hC0},
{8'hB3, 8'h85, 8'h62},
{8'hB2, 8'h70, 8'h45},
{8'hAC, 8'h57, 8'h30},
{8'hA7, 8'h49, 8'h21},
{8'hCE, 8'h84, 8'h55},
{8'hDC, 8'hB5, 8'h7B},
{8'hFB, 8'hDA, 8'hA5},
{8'hE8, 8'hAA, 8'h84},
{8'hDD, 8'h81, 8'h68},
{8'hE6, 8'h8D, 8'h60},
{8'hD4, 8'h8D, 8'h55},
{8'hCE, 8'h77, 8'h41},
{8'hE3, 8'h8F, 8'h5B},
{8'hEE, 8'hBB, 8'h84},
{8'hE6, 8'hB6, 8'h89},
{8'hD8, 8'hA8, 8'h89},
{8'hFF, 8'hF8, 8'hDB},
{8'h9D, 8'hAA, 8'h98},
{8'h51, 8'h89, 8'h73},
{8'h38, 8'h8A, 8'h71},
{8'h55, 8'h9E, 8'h86},
{8'hCE, 8'hCF, 8'hB9},
{8'hBD, 8'h80, 8'h69},
{8'hA4, 8'h50, 8'h32},
{8'hBF, 8'h7A, 8'h55},
{8'hF4, 8'hF6, 8'hC8},
{8'hFF, 8'hF6, 8'hCC},
{8'hFB, 8'hE9, 8'hBF},
{8'hD6, 8'hC1, 8'h92},
{8'hCA, 8'hA8, 8'h80},
{8'h9F, 8'h5B, 8'h41},
{8'hC0, 8'h91, 8'h78},
{8'hCF, 8'hC4, 8'hA3},
{8'hF7, 8'hF4, 8'hE4},
{8'hF4, 8'hF1, 8'hE4},
{8'hF0, 8'hEE, 8'hE2},
{8'hF4, 8'hF0, 8'hE6},
{8'hFA, 8'hF6, 8'hEC},
{8'hFB, 8'hF8, 8'hEC},
{8'hFA, 8'hF8, 8'hE8},
{8'hEF, 8'hEC, 8'hDB},
{8'hEC, 8'hEF, 8'hE3},
{8'hF5, 8'hF5, 8'hE7},
{8'hF6, 8'hF2, 8'hE1},
{8'hF2, 8'hEA, 8'hD8},
{8'hF8, 8'hF1, 8'hE0},
{8'hF5, 8'hF0, 8'hE3},
{8'hF4, 8'hF4, 8'hEB},
{8'hF9, 8'hFB, 8'hF5},
{8'hF9, 8'hF9, 8'hEF},
{8'hF7, 8'hF7, 8'hF0},
{8'hF2, 8'hF1, 8'hEE},
{8'hF4, 8'hF2, 8'hF3},
{8'hD1, 8'hCF, 8'hD2},
{8'h82, 8'h80, 8'h84},
{8'h80, 8'h7E, 8'h80},
{8'h7F, 8'h7D, 8'h7F},
{8'h7F, 8'h7D, 8'h7F},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'h7F, 8'h7D, 8'h7F},
{8'h7E, 8'h80, 8'h76},
{8'h7F, 8'h80, 8'h7B},
{8'h80, 8'h7F, 8'h83},
{8'h80, 8'h7E, 8'h89},
{8'h7B, 8'h79, 8'h86},
{8'h7B, 8'h7A, 8'h83},
{8'h7B, 8'h7B, 8'h7E},
{8'h8C, 8'h8D, 8'h87},
{8'hC7, 8'hCD, 8'hA6},
{8'hE2, 8'hE6, 8'hC6},
{8'hE7, 8'hE8, 8'hD6},
{8'hF1, 8'hF0, 8'hE7},
{8'hF2, 8'hEE, 8'hE8},
{8'hF8, 8'hF4, 8'hE9},
{8'hF9, 8'hF6, 8'hE2},
{8'hF4, 8'hF0, 8'hD2},
{8'hF3, 8'hE8, 8'hA5},
{8'hEA, 8'hEC, 8'hC3},
{8'hF0, 8'hEE, 8'hDC},
{8'hFD, 8'hEE, 8'hDC},
{8'hEB, 8'hE4, 8'hD6},
{8'hBA, 8'hC3, 8'hC3},
{8'h9D, 8'h98, 8'h94},
{8'h9E, 8'h7D, 8'h65},
{8'hAD, 8'h6C, 8'h47},
{8'hA6, 8'h52, 8'h2F},
{8'hA2, 8'h42, 8'h20},
{8'hBF, 8'h6C, 8'h44},
{8'hB4, 8'h7D, 8'h50},
{8'hDD, 8'hC1, 8'h98},
{8'hB8, 8'h8F, 8'h73},
{8'h9D, 8'h5F, 8'h4F},
{8'hE4, 8'h8D, 8'h67},
{8'hC0, 8'h7E, 8'h48},
{8'hD9, 8'h8C, 8'h59},
{8'hD9, 8'h84, 8'h51},
{8'hCC, 8'hA5, 8'h69},
{8'hFA, 8'hE1, 8'hB2},
{8'hF7, 8'hDB, 8'hBC},
{8'hFC, 8'hFF, 8'hE4},
{8'hD8, 8'hF3, 8'hD9},
{8'hA0, 8'hDF, 8'hC3},
{8'h8E, 8'hE4, 8'hCB},
{8'h83, 8'hC4, 8'hAA},
{8'hEB, 8'hF6, 8'hDA},
{8'hE1, 8'hBD, 8'h9B},
{8'hB6, 8'h68, 8'h43},
{8'hC3, 8'h7A, 8'h52},
{8'hF0, 8'hF3, 8'hC1},
{8'hFF, 8'hF4, 8'hC7},
{8'hFF, 8'hF0, 8'hC3},
{8'hBF, 8'hA8, 8'h79},
{8'hD2, 8'hAE, 8'h8A},
{8'h9E, 8'h5D, 8'h4B},
{8'hB5, 8'h86, 8'h78},
{8'hF0, 8'hEC, 8'hD8},
{8'hEE, 8'hEA, 8'hE1},
{8'hE0, 8'hDC, 8'hD3},
{8'hD9, 8'hD5, 8'hCB},
{8'hE1, 8'hDD, 8'hD2},
{8'hEE, 8'hEA, 8'hDE},
{8'hE7, 8'hE3, 8'hD5},
{8'hE9, 8'hE5, 8'hD7},
{8'hE8, 8'hE5, 8'hD6},
{8'hEA, 8'hE9, 8'hE4},
{8'hED, 8'hE9, 8'hD9},
{8'hF1, 8'hE9, 8'hC6},
{8'hF4, 8'hE9, 8'hBA},
{8'hF4, 8'hE9, 8'hB9},
{8'hED, 8'hE5, 8'hC2},
{8'hED, 8'hEA, 8'hD7},
{8'hF3, 8'hF2, 8'hEC},
{8'hF2, 8'hF1, 8'hEE},
{8'hF4, 8'hF3, 8'hF0},
{8'hFB, 8'hFA, 8'hF8},
{8'hD4, 8'hD2, 8'hD2},
{8'h8A, 8'h88, 8'h89},
{8'h7A, 8'h78, 8'h7B},
{8'hFF, 8'hD7, 8'h00},
{8'h7C, 8'h7A, 8'h7D},
{8'h7E, 8'h7C, 8'h7F},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'h7F, 8'h7D, 8'h7F},
{8'h7D, 8'h7E, 8'h78},
{8'h7E, 8'h7E, 8'h7C},
{8'h7E, 8'h7D, 8'h83},
{8'h80, 8'h7F, 8'h8A},
{8'h7F, 8'h7E, 8'h87},
{8'h7E, 8'h7E, 8'h7D},
{8'h90, 8'h92, 8'h87},
{8'hDB, 8'hDE, 8'hC9},
{8'hEC, 8'hF7, 8'hC1},
{8'hE5, 8'hF0, 8'hBD},
{8'hE3, 8'hEA, 8'hC4},
{8'hE4, 8'hE9, 8'hD0},
{8'hF2, 8'hF4, 8'hE4},
{8'hF6, 8'hF6, 8'hEB},
{8'hF8, 8'hF7, 8'hEF},
{8'hFA, 8'hF7, 8'hEC},
{8'hFB, 8'hF0, 8'hCC},
{8'hEC, 8'hEE, 8'hDE},
{8'hED, 8'hEC, 8'hE5},
{8'hFA, 8'hED, 8'hD9},
{8'hF4, 8'hF1, 8'hDF},
{8'h9D, 8'hAE, 8'hAD},
{8'h63, 8'h68, 8'h69},
{8'h7C, 8'h5C, 8'h50},
{8'h9C, 8'h59, 8'h39},
{8'hAB, 8'h5C, 8'h3C},
{8'h93, 8'h39, 8'h1A},
{8'hB7, 8'h60, 8'h40},
{8'h9D, 8'h5B, 8'h3C},
{8'h90, 8'h68, 8'h4D},
{8'h67, 8'h54, 8'h44},
{8'h2F, 8'h23, 8'h16},
{8'h96, 8'h6A, 8'h47},
{8'hE6, 8'hB7, 8'h8D},
{8'hCE, 8'h9C, 8'h6C},
{8'hE6, 8'hB6, 8'h83},
{8'hCB, 8'hA2, 8'h73},
{8'hF1, 8'hE1, 8'hBC},
{8'hFA, 8'hF5, 8'hDD},
{8'hF7, 8'hFA, 8'hE9},
{8'hEE, 8'hF8, 8'hD9},
{8'h93, 8'hAA, 8'h90},
{8'hA0, 8'hC4, 8'hB2},
{8'hC2, 8'hDC, 8'hC8},
{8'hFA, 8'hFA, 8'hDA},
{8'hEE, 8'hD3, 8'hA4},
{8'hB8, 8'h7A, 8'h49},
{8'hC2, 8'h7E, 8'h4E},
{8'hF2, 8'hF1, 8'hBD},
{8'hFF, 8'hF9, 8'hC9},
{8'hFF, 8'hF5, 8'hC5},
{8'hBC, 8'hA3, 8'h74},
{8'h90, 8'h67, 8'h45},
{8'h91, 8'h53, 8'h46},
{8'hEB, 8'hC5, 8'hC0},
{8'hF7, 8'hF8, 8'hED},
{8'hF2, 8'hF0, 8'hEA},
{8'hF2, 8'hED, 8'hE7},
{8'hED, 8'hE8, 8'hE0},
{8'hE0, 8'hDC, 8'hD1},
{8'hA3, 8'hA0, 8'h93},
{8'hB1, 8'hAE, 8'h9F},
{8'hB3, 8'hB0, 8'hA0},
{8'hE5, 8'hE2, 8'hD5},
{8'hF8, 8'hF3, 8'hF4},
{8'hF5, 8'hED, 8'hDA},
{8'hEF, 8'hE3, 8'hAD},
{8'hE9, 8'hDB, 8'h8C},
{8'hE2, 8'hD4, 8'h83},
{8'hEE, 8'hE4, 8'hA6},
{8'hF4, 8'hEE, 8'hCD},
{8'hEF, 8'hEC, 8'hE1},
{8'hF3, 8'hF1, 8'hF4},
{8'hF0, 8'hEF, 8'hF0},
{8'hBC, 8'hBB, 8'hBA},
{8'h7E, 8'h7D, 8'h7B},
{8'h7A, 8'h78, 8'h78},
{8'h7D, 8'h7B, 8'h7D},
{8'h7D, 8'h7B, 8'h7E},
{8'h7F, 8'h7D, 8'h82},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'h7F, 8'h7D, 8'h7F},
{8'h7F, 8'h7D, 8'h7F},
{8'hFF, 8'hD7, 8'h00},
{8'h7F, 8'h7D, 8'h81},
{8'h7F, 8'h7D, 8'h82},
{8'h7F, 8'h7D, 8'h82},
{8'h7F, 8'h7D, 8'h82},
{8'h7E, 8'h7D, 8'h81},
{8'h7E, 8'h7D, 8'h7D},
{8'h7D, 8'h7C, 8'h7F},
{8'h7E, 8'h7C, 8'h83},
{8'h7E, 8'h7D, 8'h83},
{8'h7E, 8'h7F, 8'h7C},
{8'h81, 8'h84, 8'h71},
{8'hD3, 8'hD9, 8'hB7},
{8'hEA, 8'hF2, 8'hC5},
{8'hDE, 8'hEE, 8'hB0},
{8'hE4, 8'hF2, 8'hB9},
{8'hE2, 8'hED, 8'hBF},
{8'hF0, 8'hF7, 8'hD7},
{8'hF8, 8'hFB, 8'hE8},
{8'hF6, 8'hF8, 8'hED},
{8'hF7, 8'hF7, 8'hF2},
{8'hF4, 8'hF3, 8'hEE},
{8'hEA, 8'hE1, 8'hCE},
{8'hEC, 8'hED, 8'hE8},
{8'hEE, 8'hEC, 8'hE9},
{8'hF5, 8'hEA, 8'hD8},
{8'hF5, 8'hF4, 8'hE2},
{8'hD7, 8'hE8, 8'hE6},
{8'h76, 8'h7C, 8'h7F},
{8'h7F, 8'h66, 8'h60},
{8'h93, 8'h50, 8'h35},
{8'hA7, 8'h58, 8'h3A},
{8'h9D, 8'h47, 8'h28},
{8'h9A, 8'h48, 8'h2A},
{8'hB6, 8'h72, 8'h58},
{8'hDD, 8'hB4, 8'hA3},
{8'h7A, 8'h79, 8'h72},
{8'h00, 8'h13, 8'h07},
{8'h35, 8'h42, 8'h21},
{8'hDE, 8'hCC, 8'hAB},
{8'hF9, 8'hEE, 8'hC3},
{8'hF1, 8'hE2, 8'hB4},
{8'hFC, 8'hD9, 8'hB5},
{8'hFC, 8'hEE, 8'hD3},
{8'hF7, 8'hFE, 8'hEC},
{8'hFD, 8'hFA, 8'hF3},
{8'hFE, 8'hF8, 8'hDA},
{8'hF7, 8'hF1, 8'hDB},
{8'hF9, 8'hF1, 8'hE5},
{8'hF9, 8'hF6, 8'hE3},
{8'hFB, 8'hF9, 8'hD3},
{8'hF1, 8'hE3, 8'hAE},
{8'hCC, 8'hA2, 8'h68},
{8'hC4, 8'h8E, 8'h57},
{8'hF2, 8'hEE, 8'hB1},
{8'hF9, 8'hEA, 8'hB9},
{8'hFF, 8'hF5, 8'hCB},
{8'hCD, 8'hAD, 8'h7E},
{8'h63, 8'h38, 8'h1B},
{8'h6E, 8'h3C, 8'h3B},
{8'hD6, 8'hB6, 8'hBF},
{8'h9F, 8'hA4, 8'hB1},
{8'hA8, 8'hA4, 8'hB4},
{8'hD6, 8'hD0, 8'hDB},
{8'hF4, 8'hF0, 8'hEC},
{8'hF2, 8'hF1, 8'hE0},
{8'hB1, 8'hB0, 8'h9D},
{8'h9F, 8'h9C, 8'h90},
{8'hD9, 8'hD7, 8'hC9},
{8'hFC, 8'hFA, 8'hE9},
{8'hFE, 8'hF8, 8'hFC},
{8'hFD, 8'hF5, 8'hE5},
{8'hF2, 8'hE7, 8'hAE},
{8'hE0, 8'hD3, 8'h7D},
{8'hE3, 8'hD7, 8'h7B},
{8'hEC, 8'hE3, 8'h9C},
{8'hF3, 8'hEC, 8'hC7},
{8'hF5, 8'hF0, 8'hE5},
{8'hF4, 8'hF2, 8'hF4},
{8'hB2, 8'hB0, 8'hB2},
{8'h74, 8'h72, 8'h72},
{8'h7D, 8'h7C, 8'h7B},
{8'h7D, 8'h7C, 8'h7A},
{8'h80, 8'h7E, 8'h7F},
{8'h83, 8'h81, 8'h85},
{8'h7F, 8'h7D, 8'h82},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'h80, 8'h7C, 8'h79},
{8'h81, 8'h7C, 8'h7B},
{8'h80, 8'h7D, 8'h81},
{8'h80, 8'h7D, 8'h85},
{8'h7F, 8'h7D, 8'h88},
{8'h7E, 8'h7D, 8'h88},
{8'h7C, 8'h7C, 8'h87},
{8'h7C, 8'h7B, 8'h85},
{8'h81, 8'h79, 8'h82},
{8'h85, 8'h7E, 8'h86},
{8'h82, 8'h7D, 8'h83},
{8'h7F, 8'h7D, 8'h7C},
{8'h75, 8'h78, 8'h69},
{8'hA4, 8'hAC, 8'h89},
{8'hE9, 8'hF5, 8'hC1},
{8'hE3, 8'hF3, 8'hB4},
{8'hE5, 8'hF1, 8'hBD},
{8'hE1, 8'hE9, 8'hC1},
{8'hE0, 8'hE3, 8'hCB},
{8'hF5, 8'hF4, 8'hE9},
{8'hF5, 8'hF2, 8'hEC},
{8'hFB, 8'hFB, 8'hEF},
{8'hED, 8'hF2, 8'hDD},
{8'hCA, 8'hD3, 8'hB5},
{8'hB5, 8'hBA, 8'h95},
{8'hC5, 8'hBE, 8'hA3},
{8'hEA, 8'hDB, 8'hCE},
{8'hF9, 8'hEA, 8'hE4},
{8'hF3, 8'hED, 8'hE7},
{8'hF7, 8'hF8, 8'hEF},
{8'h9F, 8'h9E, 8'h91},
{8'h8A, 8'h7E, 8'h6E},
{8'h8E, 8'h53, 8'h34},
{8'hA0, 8'h44, 8'h27},
{8'hAB, 8'h50, 8'h2C},
{8'h8E, 8'h51, 8'h22},
{8'hB6, 8'h87, 8'h60},
{8'hEF, 8'hCB, 8'hBD},
{8'hA3, 8'hAC, 8'hA7},
{8'h27, 8'h6A, 8'h5E},
{8'h55, 8'hAB, 8'h78},
{8'hAC, 8'hDD, 8'hB3},
{8'hF3, 8'hF9, 8'hD8},
{8'hFD, 8'hF9, 8'hD9},
{8'hFF, 8'hFD, 8'hDB},
{8'hFA, 8'hFF, 8'hE0},
{8'hFD, 8'hFB, 8'hE6},
{8'hFF, 8'hF7, 8'hE8},
{8'hF9, 8'hFA, 8'hDA},
{8'hFF, 8'hF5, 8'hDC},
{8'hFF, 8'hEF, 8'hDD},
{8'hFF, 8'hF4, 8'hDD},
{8'hFA, 8'hFA, 8'hD7},
{8'hE8, 8'hEE, 8'hBD},
{8'hCF, 8'hC5, 8'h8D},
{8'hC1, 8'hA2, 8'h69},
{8'hF6, 8'hE7, 8'h9F},
{8'hE8, 8'hE2, 8'hB1},
{8'hFC, 8'hFD, 8'hDE},
{8'hE5, 8'hA7, 8'h6D},
{8'h6C, 8'h34, 8'h2A},
{8'h1F, 8'h10, 8'h49},
{8'h7B, 8'h58, 8'h92},
{8'h56, 8'h59, 8'hAD},
{8'h5C, 8'h54, 8'hB2},
{8'h5F, 8'h52, 8'hAC},
{8'h86, 8'h7E, 8'hB4},
{8'hA0, 8'hA0, 8'h9D},
{8'hAA, 8'hAD, 8'h93},
{8'hDF, 8'hDE, 8'hD5},
{8'hF2, 8'hEF, 8'hEB},
{8'hF9, 8'hF7, 8'hE5},
{8'hF7, 8'hF0, 8'hF5},
{8'hF5, 8'hF0, 8'hF0},
{8'hEE, 8'hEA, 8'hDB},
{8'hEB, 8'hEB, 8'hC5},
{8'hED, 8'hEF, 8'hBB},
{8'hEE, 8'hEF, 8'hC2},
{8'hF2, 8'hEF, 8'hDD},
{8'hFA, 8'hF4, 8'hF7},
{8'hFC, 8'hFB, 8'hF9},
{8'hEC, 8'hEB, 8'hE8},
{8'h96, 8'h95, 8'h93},
{8'h79, 8'h78, 8'h77},
{8'h7E, 8'h7C, 8'h7E},
{8'h81, 8'h7F, 8'h82},
{8'h7E, 8'h7C, 8'h80},
{8'h7E, 8'h7C, 8'h81},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'h81, 8'h7C, 8'h7F},
{8'h80, 8'h7D, 8'h80},
{8'h80, 8'h7E, 8'h81},
{8'h80, 8'h7F, 8'h82},
{8'h7E, 8'h7E, 8'h80},
{8'h7F, 8'h80, 8'h82},
{8'h7D, 8'h7F, 8'h7F},
{8'h78, 8'h7A, 8'h7B},
{8'h80, 8'h7A, 8'h81},
{8'h81, 8'h7B, 8'h83},
{8'h80, 8'h7B, 8'h85},
{8'h80, 8'h7E, 8'h83},
{8'h7D, 8'h7E, 8'h78},
{8'hCE, 8'hD3, 8'hBE},
{8'hEE, 8'hF8, 8'hD1},
{8'hE5, 8'hF1, 8'hC2},
{8'hD7, 8'hE3, 8'hB5},
{8'hA9, 8'hB0, 8'h8D},
{8'hE1, 8'hE3, 8'hCF},
{8'hF5, 8'hF2, 8'hE9},
{8'hF3, 8'hF0, 8'hE9},
{8'hE6, 8'hE8, 8'hD9},
{8'hE5, 8'hEA, 8'hD1},
{8'hC7, 8'hD1, 8'hAE},
{8'hC3, 8'hCA, 8'h9C},
{8'hB8, 8'hB2, 8'h8E},
{8'hB4, 8'hA5, 8'h91},
{8'hF8, 8'hEC, 8'hE2},
{8'hEE, 8'hE9, 8'hE1},
{8'hF5, 8'hF5, 8'hED},
{8'h9D, 8'h98, 8'h8E},
{8'h84, 8'h74, 8'h67},
{8'hA9, 8'h6F, 8'h4B},
{8'hAD, 8'h57, 8'h35},
{8'hAD, 8'h54, 8'h31},
{8'h97, 8'h52, 8'h2B},
{8'h8E, 8'h53, 8'h34},
{8'hF7, 8'hD6, 8'hC6},
{8'hF3, 8'hF2, 8'hE8},
{8'h9C, 8'hD2, 8'hBE},
{8'hA9, 8'hDD, 8'hB5},
{8'hBB, 8'hD3, 8'hAE},
{8'hFA, 8'hF8, 8'hDA},
{8'hF3, 8'hE8, 8'hC9},
{8'hFF, 8'hFF, 8'hDD},
{8'hF8, 8'hFF, 8'hDE},
{8'hF8, 8'hFF, 8'hE3},
{8'hFA, 8'hFD, 8'hE6},
{8'hF4, 8'hFF, 8'hDA},
{8'hFC, 8'hFA, 8'hDC},
{8'hFF, 8'hF5, 8'hDF},
{8'hFF, 8'hF8, 8'hE1},
{8'hFB, 8'hFC, 8'hDD},
{8'hEF, 8'hED, 8'hC5},
{8'hF3, 8'hDF, 8'hB2},
{8'hDB, 8'hAE, 8'h85},
{8'hEF, 8'hE5, 8'hBB},
{8'hDC, 8'hCF, 8'h89},
{8'hF9, 8'hFE, 8'hC4},
{8'hD0, 8'hA5, 8'h67},
{8'h84, 8'h40, 8'h34},
{8'h51, 8'h3A, 8'h80},
{8'h81, 8'h76, 8'hB7},
{8'h7D, 8'h7E, 8'hAD},
{8'h6A, 8'h5E, 8'hB0},
{8'h6A, 8'h5C, 8'hAE},
{8'h5C, 8'h4D, 8'hA1},
{8'h5D, 8'h4E, 8'h98},
{8'h81, 8'h76, 8'h9D},
{8'hD7, 8'hD1, 8'hD4},
{8'hF2, 8'hEC, 8'hE7},
{8'hF7, 8'hEF, 8'hF6},
{8'hFD, 8'hF9, 8'hF3},
{8'hF5, 8'hF0, 8'hE9},
{8'hF2, 8'hEE, 8'hE3},
{8'hFB, 8'hFA, 8'hE1},
{8'hE9, 8'hE9, 8'hC5},
{8'hEF, 8'hEF, 8'hCE},
{8'hF8, 8'hF4, 8'hE9},
{8'hFA, 8'hF4, 8'hF9},
{8'hF8, 8'hF7, 8'hF4},
{8'hFD, 8'hFC, 8'hF9},
{8'hE0, 8'hDF, 8'hDD},
{8'h86, 8'h85, 8'h84},
{8'h7D, 8'h7B, 8'h7D},
{8'h85, 8'h83, 8'h86},
{8'h7C, 8'h7A, 8'h7E},
{8'h7F, 8'h7D, 8'h82},
{8'h80, 8'h7E, 8'h81},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'h80, 8'h7C, 8'h85},
{8'h80, 8'h7D, 8'h85},
{8'h80, 8'h7F, 8'h81},
{8'h7F, 8'h80, 8'h7D},
{8'h7A, 8'h7C, 8'h73},
{8'h75, 8'h7A, 8'h6D},
{8'h78, 8'h7F, 8'h6F},
{8'h80, 8'h87, 8'h77},
{8'h87, 8'h85, 8'h80},
{8'h8E, 8'h8C, 8'h8B},
{8'h8A, 8'h89, 8'h8B},
{8'h79, 8'h7A, 8'h7C},
{8'h7A, 8'h7C, 8'h79},
{8'hB3, 8'hB7, 8'hA9},
{8'hC8, 8'hD0, 8'hB6},
{8'hC6, 8'hD1, 8'hAD},
{8'hBB, 8'hC5, 8'h9F},
{8'hC6, 8'hCC, 8'hAF},
{8'hF2, 8'hF3, 8'hE3},
{8'hE8, 8'hE5, 8'hDD},
{8'hB5, 8'hB3, 8'hAB},
{8'hB2, 8'hB4, 8'hA2},
{8'hF0, 8'hF6, 8'hD9},
{8'hDE, 8'hE9, 8'hC1},
{8'hCB, 8'hD5, 8'h9C},
{8'hBA, 8'hB9, 8'h8B},
{8'hA8, 8'h9B, 8'h7E},
{8'hCC, 8'hC0, 8'hB0},
{8'hF1, 8'hED, 8'hE3},
{8'hE9, 8'hE7, 8'hDF},
{8'h98, 8'h8C, 8'h86},
{8'h7E, 8'h66, 8'h5D},
{8'hBF, 8'h92, 8'h66},
{8'hC1, 8'h78, 8'h50},
{8'hB7, 8'h63, 8'h43},
{8'h8F, 8'h40, 8'h24},
{8'h90, 8'h43, 8'h2E},
{8'hCB, 8'h90, 8'h80},
{8'hFF, 8'hF8, 8'hE1},
{8'hBE, 8'hDA, 8'hB7},
{8'h99, 8'hA9, 8'h88},
{8'hE7, 8'hE4, 8'hC8},
{8'hFE, 8'hF7, 8'hDD},
{8'hF0, 8'hE2, 8'hC5},
{8'hFE, 8'hFC, 8'hDB},
{8'hFB, 8'hFF, 8'hDE},
{8'hFA, 8'hFF, 8'hE1},
{8'hFB, 8'hFF, 8'hE4},
{8'hF9, 8'hFF, 8'hDA},
{8'hFD, 8'hFF, 8'hDD},
{8'hFF, 8'hFB, 8'hE0},
{8'hFF, 8'hFC, 8'hE4},
{8'hFB, 8'hF9, 8'hDF},
{8'hF1, 8'hEC, 8'hCD},
{8'hFF, 8'hEB, 8'hCB},
{8'hE3, 8'hB1, 8'h91},
{8'hEA, 8'hDF, 8'hB6},
{8'hD8, 8'hCA, 8'h7E},
{8'hFE, 8'hFF, 8'hCC},
{8'hBF, 8'h9D, 8'h6F},
{8'h99, 8'h4D, 8'h31},
{8'h52, 8'h37, 8'h58},
{8'h45, 8'h48, 8'h7E},
{8'h63, 8'h58, 8'h83},
{8'h43, 8'h33, 8'h7B},
{8'h30, 8'h25, 8'h4C},
{8'h23, 8'h1A, 8'h3C},
{8'h1C, 8'h0D, 8'h56},
{8'h3A, 8'h25, 8'h77},
{8'h84, 8'h76, 8'h92},
{8'hF8, 8'hF3, 8'hE1},
{8'hFC, 8'hF7, 8'hDA},
{8'hF0, 8'hEE, 8'hD5},
{8'hF4, 8'hF0, 8'hE2},
{8'hF8, 8'hF3, 8'hED},
{8'hF7, 8'hF2, 8'hEA},
{8'hF6, 8'hF4, 8'hE4},
{8'hE3, 8'hE1, 8'hD1},
{8'hF6, 8'hF2, 8'hED},
{8'hFD, 8'hF8, 8'hFC},
{8'hFB, 8'hFA, 8'hF6},
{8'hF8, 8'hF7, 8'hF4},
{8'hFC, 8'hFC, 8'hFA},
{8'hC2, 8'hC1, 8'hC0},
{8'h7C, 8'h7A, 8'h7C},
{8'h82, 8'h80, 8'h83},
{8'h84, 8'h82, 8'h86},
{8'h7F, 8'h7D, 8'h82},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'h7F, 8'h7D, 8'h81},
{8'h80, 8'h7C, 8'h8A},
{8'h80, 8'h7F, 8'h88},
{8'h80, 8'h81, 8'h80},
{8'h8B, 8'h8E, 8'h82},
{8'hA3, 8'hAA, 8'h93},
{8'h91, 8'h9A, 8'h7D},
{8'hA3, 8'hAE, 8'h8C},
{8'hCD, 8'hD8, 8'hB7},
{8'hD6, 8'hDC, 8'hBE},
{8'hDD, 8'hE2, 8'hC9},
{8'hA0, 8'hA4, 8'h92},
{8'h7D, 8'h80, 8'h73},
{8'h79, 8'h7C, 8'h6F},
{8'h74, 8'h79, 8'h64},
{8'h94, 8'h9B, 8'h7E},
{8'hDD, 8'hE5, 8'hC2},
{8'hC1, 8'hCB, 8'hA9},
{8'hC4, 8'hCA, 8'hB2},
{8'hD3, 8'hD4, 8'hC8},
{8'hAB, 8'hA9, 8'hA3},
{8'hE6, 8'hE4, 8'hDD},
{8'h90, 8'h92, 8'h81},
{8'hBD, 8'hC3, 8'hA4},
{8'hE8, 8'hF4, 8'hC9},
{8'hD1, 8'hDB, 8'hA0},
{8'hAC, 8'hAD, 8'h7C},
{8'hB2, 8'hA9, 8'h88},
{8'hB1, 8'hA9, 8'h95},
{8'hBD, 8'hBB, 8'hAE},
{8'hD7, 8'hD3, 8'hC9},
{8'h9D, 8'h8B, 8'h85},
{8'h79, 8'h58, 8'h4F},
{8'hC5, 8'hA6, 8'h73},
{8'hC8, 8'h92, 8'h63},
{8'hBA, 8'h6F, 8'h4E},
{8'h89, 8'h32, 8'h1D},
{8'h9F, 8'h45, 8'h37},
{8'h95, 8'h4E, 8'h3D},
{8'hF4, 8'hDC, 8'hBC},
{8'hF3, 8'hF8, 8'hCF},
{8'hF6, 8'hF7, 8'hD7},
{8'hFF, 8'hF9, 8'hDC},
{8'hFB, 8'hF3, 8'hD7},
{8'hFF, 8'hF8, 8'hDB},
{8'hFF, 8'hFB, 8'hDC},
{8'hFF, 8'hFE, 8'hDF},
{8'hFB, 8'hF4, 8'hD6},
{8'hF6, 8'hEE, 8'hCF},
{8'hFA, 8'hEF, 8'hCD},
{8'hF9, 8'hF1, 8'hD2},
{8'hFF, 8'hFC, 8'hE1},
{8'hFF, 8'hFE, 8'hE6},
{8'hF5, 8'hF3, 8'hD9},
{8'hF5, 8'hEF, 8'hD3},
{8'hFC, 8'hE9, 8'hCB},
{8'hDC, 8'hB3, 8'h91},
{8'hD6, 8'hC4, 8'h86},
{8'hD9, 8'hC9, 8'h90},
{8'hFF, 8'hF6, 8'hD9},
{8'hB5, 8'h7F, 8'h66},
{8'h9C, 8'h52, 8'h2A},
{8'h41, 8'h20, 8'h10},
{8'h23, 8'h1B, 8'h38},
{8'h22, 8'h13, 8'h4B},
{8'h25, 8'h1E, 8'h28},
{8'h07, 8'h00, 8'h0A},
{8'h1E, 8'h16, 8'h2E},
{8'h3B, 8'h30, 8'h51},
{8'h83, 8'h78, 8'h83},
{8'hCF, 8'hC9, 8'hAD},
{8'hD8, 8'hD6, 8'hAC},
{8'hC2, 8'hBB, 8'h99},
{8'hC8, 8'hC7, 8'hA6},
{8'hF9, 8'hF7, 8'hE7},
{8'hF6, 8'hF0, 8'hF0},
{8'hF7, 8'hF0, 8'hF6},
{8'hFA, 8'hF6, 8'hF4},
{8'hA5, 8'hA1, 8'h9A},
{8'h95, 8'h8F, 8'h8C},
{8'hDB, 8'hD6, 8'hD9},
{8'hF0, 8'hEF, 8'hEB},
{8'hFA, 8'hFA, 8'hF7},
{8'hFD, 8'hFD, 8'hFB},
{8'hF5, 8'hF3, 8'hF3},
{8'h9A, 8'h98, 8'h9A},
{8'h77, 8'h75, 8'h78},
{8'h7D, 8'h7B, 8'h7F},
{8'h7C, 8'h7A, 8'h7F},
{8'h7E, 8'h7C, 8'h7F},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'h7E, 8'h7C, 8'h81},
{8'h7E, 8'h7C, 8'h8B},
{8'h7D, 8'h7D, 8'h85},
{8'h76, 8'h78, 8'h70},
{8'hA8, 8'hAF, 8'h97},
{8'hEA, 8'hF4, 8'hD0},
{8'hE4, 8'hF1, 8'hC5},
{8'hE3, 8'hF1, 8'hC2},
{8'hE4, 8'hF2, 8'hC1},
{8'hE3, 8'hF1, 8'hBA},
{8'hC4, 8'hD1, 8'h9E},
{8'hCE, 8'hD9, 8'hB0},
{8'hD2, 8'hDB, 8'hBA},
{8'hB8, 8'hC0, 8'hA1},
{8'hB3, 8'hBB, 8'h99},
{8'hC5, 8'hCD, 8'hA3},
{8'hB2, 8'hBB, 8'h8E},
{8'hC9, 8'hD2, 8'hB1},
{8'hD0, 8'hD4, 8'hBD},
{8'h81, 8'h82, 8'h76},
{8'hBA, 8'hB7, 8'hB3},
{8'hFD, 8'hF9, 8'hF5},
{8'hC0, 8'hC1, 8'hB2},
{8'h91, 8'h97, 8'h7A},
{8'hDA, 8'hE5, 8'hBC},
{8'hE7, 8'hF0, 8'hBD},
{8'hBC, 8'hBD, 8'h93},
{8'hA7, 8'hA0, 8'h84},
{8'hCC, 8'hC5, 8'hB3},
{8'h8C, 8'h8A, 8'h7B},
{8'h98, 8'h92, 8'h84},
{8'h93, 8'h7B, 8'h70},
{8'h7F, 8'h57, 8'h49},
{8'hCD, 8'hAD, 8'h7A},
{8'hD9, 8'hB3, 8'h81},
{8'hBC, 8'h7F, 8'h59},
{8'h8F, 8'h35, 8'h20},
{8'h9D, 8'h3C, 8'h2D},
{8'h8A, 8'h43, 8'h2F},
{8'hC0, 8'hA1, 8'h80},
{8'hFF, 8'hFD, 8'hD6},
{8'hFA, 8'hF9, 8'hD8},
{8'hF8, 8'hFB, 8'hDA},
{8'hFB, 8'hFB, 8'hDB},
{8'hFE, 8'hFE, 8'hDF},
{8'hF5, 8'hE7, 8'hCA},
{8'hEA, 8'hCB, 8'hB2},
{8'hEF, 8'hC3, 8'hA9},
{8'hEE, 8'hBC, 8'hA2},
{8'hF4, 8'hBC, 8'hA6},
{8'hE2, 8'hBE, 8'hA5},
{8'hFC, 8'hF7, 8'hDD},
{8'hFD, 8'hFD, 8'hE3},
{8'hEA, 8'hE9, 8'hCD},
{8'hFC, 8'hF8, 8'hD8},
{8'hF4, 8'hE6, 8'hC3},
{8'hD9, 8'hB8, 8'h8E},
{8'hD2, 8'hA4, 8'h69},
{8'hE1, 8'hD7, 8'hAF},
{8'hFC, 8'hE1, 8'hBA},
{8'hAD, 8'h5C, 8'h41},
{8'h84, 8'h41, 8'h2D},
{8'h64, 8'h3B, 8'h20},
{8'h2A, 8'h11, 8'h1D},
{8'h1A, 8'h0D, 8'h49},
{8'h26, 8'h20, 8'h30},
{8'h1C, 8'h14, 8'h2A},
{8'h8B, 8'h82, 8'h8C},
{8'hE3, 8'hDF, 8'hC5},
{8'hF6, 8'hF4, 8'hD0},
{8'hDA, 8'hD3, 8'hBF},
{8'hAE, 8'hA5, 8'h93},
{8'hAD, 8'hA7, 8'h82},
{8'hC1, 8'hC0, 8'hA3},
{8'hFA, 8'hF8, 8'hEE},
{8'hF9, 8'hF3, 8'hF8},
{8'hF8, 8'hF0, 8'hFA},
{8'hF3, 8'hEE, 8'hEE},
{8'h90, 8'h8C, 8'h83},
{8'h76, 8'h71, 8'h68},
{8'hD7, 8'hD3, 8'hCF},
{8'hD3, 8'hD2, 8'hCE},
{8'h94, 8'h93, 8'h90},
{8'hC6, 8'hC6, 8'hC3},
{8'hDE, 8'hDC, 8'hDC},
{8'h91, 8'h8F, 8'h91},
{8'h7A, 8'h78, 8'h7B},
{8'h80, 8'h7E, 8'h82},
{8'h7E, 8'h7C, 8'h81},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'h7F, 8'h7D, 8'h81},
{8'h7B, 8'h7B, 8'h86},
{8'h78, 8'h79, 8'h7B},
{8'h78, 8'h7D, 8'h6D},
{8'h9D, 8'hA7, 8'h84},
{8'hE5, 8'hF2, 8'hC2},
{8'hE3, 8'hF2, 8'hBC},
{8'hE0, 8'hF1, 8'hBA},
{8'hDF, 8'hF0, 8'hB7},
{8'hDE, 8'hF2, 8'hAE},
{8'hDE, 8'hF1, 8'hB3},
{8'hE6, 8'hF6, 8'hC1},
{8'hE6, 8'hF3, 8'hC7},
{8'hE8, 8'hF3, 8'hCB},
{8'hE8, 8'hF1, 8'hC7},
{8'hE3, 8'hEC, 8'hBC},
{8'hD4, 8'hDD, 8'hAA},
{8'hBF, 8'hC9, 8'hA4},
{8'h81, 8'h86, 8'h6B},
{8'h7C, 8'h7D, 8'h70},
{8'hE3, 8'hE0, 8'hDC},
{8'hF8, 8'hF5, 8'hF2},
{8'hF0, 8'hF1, 8'hE5},
{8'hD6, 8'hDB, 8'hC3},
{8'h9B, 8'hA5, 8'h83},
{8'hCC, 8'hD3, 8'hB4},
{8'hA5, 8'hA4, 8'h8D},
{8'hAF, 8'hA8, 8'h98},
{8'hBC, 8'hB6, 8'hAA},
{8'hAD, 8'hAB, 8'h9C},
{8'h8E, 8'h86, 8'h72},
{8'h9E, 8'h82, 8'h6C},
{8'h8F, 8'h60, 8'h49},
{8'hBE, 8'hA2, 8'h73},
{8'hEB, 8'hDA, 8'hA5},
{8'hC0, 8'h93, 8'h64},
{8'h96, 8'h3F, 8'h21},
{8'h96, 8'h35, 8'h20},
{8'h92, 8'h53, 8'h3C},
{8'h90, 8'h75, 8'h5A},
{8'hEC, 8'hE1, 8'hC7},
{8'hFF, 8'hFF, 8'hDE},
{8'hF9, 8'hFE, 8'hDB},
{8'hF6, 8'hFF, 8'hDF},
{8'hFE, 8'hFF, 8'hE2},
{8'hE7, 8'hCF, 8'hB2},
{8'hE5, 8'hAF, 8'h97},
{8'hFE, 8'hC1, 8'hA8},
{8'hFE, 8'hBE, 8'hA2},
{8'hFF, 8'hBE, 8'hAD},
{8'hED, 8'hC1, 8'hAB},
{8'hFB, 8'hF7, 8'hDB},
{8'hF9, 8'hFA, 8'hDC},
{8'hEB, 8'hE5, 8'hC6},
{8'hFF, 8'hF9, 8'hD7},
{8'hDA, 8'hBE, 8'h96},
{8'hCB, 8'hA1, 8'h73},
{8'hC9, 8'h88, 8'h62},
{8'hF5, 8'hF0, 8'hC8},
{8'hE3, 8'hBA, 8'h71},
{8'hA4, 8'h53, 8'h2E},
{8'h66, 8'h2E, 8'h2F},
{8'h6A, 8'h43, 8'h2E},
{8'h19, 8'h0C, 8'h11},
{8'h09, 8'h05, 8'h38},
{8'h2D, 8'h22, 8'h5B},
{8'h19, 8'h0D, 8'h41},
{8'h3D, 8'h37, 8'h45},
{8'hCB, 8'hCB, 8'hA9},
{8'hD5, 8'hD4, 8'hB6},
{8'hFB, 8'hF4, 8'hF8},
{8'hE6, 8'hDC, 8'hE6},
{8'hC3, 8'hBB, 8'hAC},
{8'hC7, 8'hC3, 8'hBA},
{8'hFF, 8'hFA, 8'hFE},
{8'hFF, 8'hFA, 8'hFF},
{8'hFB, 8'hF6, 8'hFA},
{8'hF3, 8'hF1, 8'hE5},
{8'hBE, 8'hBC, 8'hA6},
{8'hB2, 8'hAF, 8'h9B},
{8'hEC, 8'hE9, 8'hDB},
{8'hEE, 8'hED, 8'hE8},
{8'h8F, 8'h8E, 8'h8B},
{8'h75, 8'h74, 8'h72},
{8'h7F, 8'h7E, 8'h7D},
{8'h7B, 8'h79, 8'h7B},
{8'hFF, 8'hD7, 8'h00},
{8'h7D, 8'h7B, 8'h7F},
{8'h7D, 8'h7B, 8'h80},
{8'h7F, 8'h7D, 8'h81},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'h7D, 8'h7E, 8'h85},
{8'h7A, 8'h7D, 8'h79},
{8'h91, 8'h99, 8'h83},
{8'hC6, 8'hD2, 8'hA8},
{8'hE5, 8'hF3, 8'hBC},
{8'hE1, 8'hF3, 8'hB6},
{8'hE0, 8'hF2, 8'hB6},
{8'hDE, 8'hF2, 8'hB6},
{8'hDC, 8'hF1, 8'hB1},
{8'hE3, 8'hF6, 8'hBD},
{8'hE1, 8'hF2, 8'hC1},
{8'hD0, 8'hDE, 8'hB6},
{8'hDA, 8'hE4, 8'hC0},
{8'hE3, 8'hEC, 8'hC4},
{8'hE1, 8'hE9, 8'hBC},
{8'hEC, 8'hF4, 8'hC3},
{8'hC4, 8'hCF, 8'hA6},
{8'h8A, 8'h90, 8'h72},
{8'h91, 8'h92, 8'h83},
{8'hF7, 8'hF5, 8'hF1},
{8'hF5, 8'hF1, 8'hF0},
{8'hF3, 8'hF3, 8'hED},
{8'hD7, 8'hDB, 8'hCA},
{8'h74, 8'h7C, 8'h64},
{8'h83, 8'h88, 8'h7D},
{8'hB2, 8'hB1, 8'hAC},
{8'hEB, 8'hE5, 8'hE3},
{8'hEC, 8'hE8, 8'hE3},
{8'hF5, 8'hF5, 8'hE8},
{8'hCC, 8'hC2, 8'hAB},
{8'hD2, 8'hB9, 8'h99},
{8'h91, 8'h62, 8'h3F},
{8'hA0, 8'h82, 8'h57},
{8'hFE, 8'hFC, 8'hC6},
{8'hD5, 8'hB7, 8'h7F},
{8'hA9, 8'h58, 8'h30},
{8'h99, 8'h3C, 8'h20},
{8'h72, 8'h3F, 8'h24},
{8'h7E, 8'h6B, 8'h5A},
{8'h9E, 8'h8A, 8'h83},
{8'hF5, 8'hE1, 8'hC6},
{8'hFF, 8'hFF, 8'hDE},
{8'hF7, 8'hFF, 8'hE1},
{8'hF9, 8'hFF, 8'hDF},
{8'hFC, 8'hEE, 8'hD0},
{8'hEF, 8'hBB, 8'hA1},
{8'hFC, 8'hBC, 8'h9E},
{8'hFE, 8'hC0, 8'h9C},
{8'hFB, 8'hB9, 8'hA7},
{8'hF4, 8'hD1, 8'hB8},
{8'hFF, 8'hFE, 8'hDF},
{8'hF6, 8'hF9, 8'hD9},
{8'hF1, 8'hE6, 8'hC5},
{8'hFB, 8'hDA, 8'hB8},
{8'hBF, 8'h80, 8'h57},
{8'hD6, 8'h94, 8'h65},
{8'hCD, 8'h99, 8'h6D},
{8'hF9, 8'hF4, 8'hBB},
{8'hB1, 8'h88, 8'h40},
{8'h8E, 8'h54, 8'h3F},
{8'hBC, 8'h8E, 8'h7C},
{8'h86, 8'h70, 8'h41},
{8'h2D, 8'h4F, 8'h59},
{8'h57, 8'h61, 8'h97},
{8'h8C, 8'h83, 8'hB0},
{8'h80, 8'h78, 8'hA2},
{8'h5E, 8'h57, 8'h7D},
{8'h9D, 8'h98, 8'hA3},
{8'hCE, 8'hCC, 8'hBA},
{8'hF9, 8'hF8, 8'hDF},
{8'hFB, 8'hF8, 8'hF1},
{8'hF1, 8'hE8, 8'hF8},
{8'hA8, 8'hA0, 8'hAF},
{8'hA6, 8'h9F, 8'hAC},
{8'hDA, 8'hD3, 8'hDE},
{8'hFD, 8'hFA, 8'hF5},
{8'hF5, 8'hF3, 8'hDA},
{8'hF4, 8'hF5, 8'hD0},
{8'hE6, 8'hE6, 8'hC5},
{8'hEC, 8'hEA, 8'hD4},
{8'hED, 8'hEC, 8'hE7},
{8'h9B, 8'h9A, 8'h98},
{8'h79, 8'h77, 8'h76},
{8'h83, 8'h81, 8'h81},
{8'h81, 8'h7F, 8'h81},
{8'h7E, 8'h7C, 8'h7F},
{8'h7E, 8'h7C, 8'h80},
{8'h7D, 8'h7B, 8'h80},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'h7F, 8'h7D, 8'h7F},
{8'h7F, 8'h7D, 8'h7F},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'h7F, 8'h7D, 8'h7F},
{8'hFF, 8'hD7, 8'h00},
{8'h76, 8'h78, 8'h7A},
{8'hA1, 8'hA7, 8'h98},
{8'hE5, 8'hEF, 8'hCD},
{8'hE7, 8'hF4, 8'hC5},
{8'hE3, 8'hF3, 8'hBB},
{8'hE1, 8'hF4, 8'hB4},
{8'hE0, 8'hF3, 8'hB5},
{8'hDE, 8'hF2, 8'hB7},
{8'hDF, 8'hF5, 8'hB7},
{8'hE1, 8'hF3, 8'hBD},
{8'hD9, 8'hE8, 8'hBF},
{8'hD5, 8'hDF, 8'hC0},
{8'hF2, 8'hF8, 8'hDF},
{8'hE3, 8'hE8, 8'hCC},
{8'hE4, 8'hEA, 8'hC7},
{8'hE5, 8'hEC, 8'hC2},
{8'hE3, 8'hF0, 8'hBB},
{8'hB5, 8'hBE, 8'h93},
{8'hBC, 8'hBF, 8'hA7},
{8'hFF, 8'hFC, 8'hF4},
{8'hF4, 8'hF0, 8'hF0},
{8'hF2, 8'hF2, 8'hEB},
{8'hCF, 8'hD3, 8'hBE},
{8'hA7, 8'hAE, 8'h91},
{8'hE6, 8'hE4, 8'hE7},
{8'hFD, 8'hF9, 8'hFE},
{8'hFC, 8'hF7, 8'hF7},
{8'hF7, 8'hF3, 8'hEF},
{8'hFB, 8'hF9, 8'hEE},
{8'hD6, 8'hCA, 8'hAD},
{8'hE2, 8'hC7, 8'hA2},
{8'h8C, 8'h5B, 8'h3E},
{8'h93, 8'h77, 8'h5B},
{8'hF6, 8'hF6, 8'hC7},
{8'hF5, 8'hE3, 8'hA7},
{8'hCD, 8'h85, 8'h51},
{8'h97, 8'h43, 8'h1B},
{8'h6A, 8'h38, 8'h1A},
{8'h7D, 8'h67, 8'h58},
{8'h87, 8'h71, 8'h6F},
{8'hA4, 8'h7A, 8'h6A},
{8'hE0, 8'hD1, 8'hB1},
{8'hF7, 8'hFD, 8'hDA},
{8'hF7, 8'hFF, 8'hDE},
{8'hFE, 8'hF9, 8'hDA},
{8'hFB, 8'hDE, 8'hBF},
{8'hFA, 8'hCD, 8'hAA},
{8'hF7, 8'hC8, 8'hAA},
{8'hF9, 8'hC7, 8'hB4},
{8'hFA, 8'hEC, 8'hCD},
{8'hF7, 8'hFF, 8'hDE},
{8'hEB, 8'hF4, 8'hCE},
{8'hF2, 8'hDA, 8'hB8},
{8'hD0, 8'h8A, 8'h6D},
{8'hC2, 8'h6B, 8'h47},
{8'hC8, 8'h71, 8'h43},
{8'hDE, 8'hB8, 8'h7F},
{8'hC6, 8'hB4, 8'h87},
{8'h66, 8'h53, 8'h41},
{8'h4F, 8'h47, 8'h5D},
{8'hBB, 8'h9F, 8'h7F},
{8'hDF, 8'hD6, 8'h7C},
{8'h44, 8'h75, 8'h6D},
{8'h3A, 8'h4F, 8'h98},
{8'h62, 8'h60, 8'hAC},
{8'hA0, 8'hA4, 8'hC2},
{8'hAE, 8'hB5, 8'hBD},
{8'h8A, 8'h8E, 8'h97},
{8'hC8, 8'hCB, 8'hC8},
{8'hF9, 8'hFC, 8'hE6},
{8'hFF, 8'hFE, 8'hEA},
{8'hB9, 8'hB5, 8'hB9},
{8'h1F, 8'h18, 8'h30},
{8'h05, 8'h00, 8'h18},
{8'h1E, 8'h14, 8'h24},
{8'h52, 8'h4C, 8'h40},
{8'hC2, 8'hC0, 8'h91},
{8'hF1, 8'hF1, 8'hBB},
{8'hE8, 8'hE8, 8'hBB},
{8'hEA, 8'hE9, 8'hC7},
{8'hE8, 8'hE7, 8'hDF},
{8'h9D, 8'h9C, 8'h98},
{8'h79, 8'h79, 8'h75},
{8'hB0, 8'hAF, 8'hAE},
{8'h96, 8'h94, 8'h97},
{8'h7A, 8'h78, 8'h7C},
{8'h80, 8'h7E, 8'h82},
{8'h7F, 8'h7D, 8'h81},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'h7F, 8'h7E, 8'h7B},
{8'h7F, 8'h7E, 8'h7C},
{8'h7F, 8'h7D, 8'h7E},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'h7F, 8'h7D, 8'h7E},
{8'h7F, 8'h7E, 8'h7C},
{8'h7E, 8'h7D, 8'h7B},
{8'h7B, 8'h7F, 8'h7C},
{8'hCB, 8'hD8, 8'hAB},
{8'hE6, 8'hF7, 8'hB4},
{8'hDE, 8'hEE, 8'hBB},
{8'hE0, 8'hF1, 8'hC2},
{8'hE1, 8'hF6, 8'hB5},
{8'hE0, 8'hF6, 8'hB3},
{8'hE0, 8'hF4, 8'hC0},
{8'hDF, 8'hF4, 8'hAB},
{8'hE7, 8'hF5, 8'hB9},
{8'hE4, 8'hEC, 8'hC6},
{8'hF2, 8'hF1, 8'hE1},
{8'hF4, 8'hF1, 8'hEA},
{8'hF1, 8'hF0, 8'hE7},
{8'hEA, 8'hEC, 8'hDD},
{8'hE5, 8'hEB, 8'hD2},
{8'hE2, 8'hF2, 8'hBF},
{8'hDD, 8'hE9, 8'hB8},
{8'hD5, 8'hD9, 8'hB6},
{8'hF9, 8'hF8, 8'hE8},
{8'hFA, 8'hF4, 8'hF4},
{8'hF9, 8'hF5, 8'hF3},
{8'hE6, 8'hE8, 8'hD2},
{8'hF9, 8'hFB, 8'hDB},
{8'hFF, 8'hF6, 8'hFF},
{8'hFD, 8'hF2, 8'hF8},
{8'hF9, 8'hF8, 8'hE6},
{8'hF9, 8'hF6, 8'hEF},
{8'hFF, 8'hF8, 8'hFF},
{8'hC7, 8'hB7, 8'h95},
{8'hE2, 8'hCE, 8'h98},
{8'h9D, 8'h74, 8'h72},
{8'hB1, 8'h91, 8'h90},
{8'hD0, 8'hB5, 8'h98},
{8'hFF, 8'hFE, 8'hBD},
{8'hE3, 8'hC3, 8'h76},
{8'h9E, 8'h51, 8'h20},
{8'h74, 8'h30, 8'h1C},
{8'h8C, 8'h75, 8'h6C},
{8'h83, 8'h7A, 8'h7C},
{8'h96, 8'h81, 8'h7D},
{8'hD5, 8'hC8, 8'hA0},
{8'hD2, 8'hCA, 8'h9B},
{8'hF2, 8'hEE, 8'hDA},
{8'hFF, 8'hFF, 8'hEE},
{8'hFF, 8'hFF, 8'hD6},
{8'hF9, 8'hF6, 8'hD3},
{8'hF6, 8'hEC, 8'hEB},
{8'hFC, 8'hF4, 8'hE5},
{8'hFA, 8'hFE, 8'hDC},
{8'hF6, 8'hFF, 8'hD6},
{8'hEC, 8'hE2, 8'hB5},
{8'hC8, 8'h87, 8'h6D},
{8'hB5, 8'h53, 8'h41},
{8'hC4, 8'h6A, 8'h49},
{8'hBD, 8'h78, 8'h43},
{8'hE7, 8'hBC, 8'h97},
{8'h64, 8'h4D, 8'h7B},
{8'h17, 8'h4B, 8'hAC},
{8'h03, 8'h60, 8'hBD},
{8'h39, 8'h5E, 8'h7D},
{8'hE4, 8'hBE, 8'h76},
{8'hD2, 8'hB8, 8'h77},
{8'h31, 8'h55, 8'h88},
{8'h16, 8'h3B, 8'h92},
{8'h22, 8'h42, 8'h97},
{8'h38, 8'h54, 8'h96},
{8'h70, 8'h88, 8'hA3},
{8'hA0, 8'hB4, 8'hA9},
{8'hC8, 8'hD5, 8'hBF},
{8'h95, 8'h97, 8'h93},
{8'h22, 8'h1F, 8'h30},
{8'h00, 8'h03, 8'h12},
{8'h0C, 8'h07, 8'h2C},
{8'h36, 8'h28, 8'h3A},
{8'h97, 8'h89, 8'h5B},
{8'hDE, 8'hD2, 8'h77},
{8'hF3, 8'hE8, 8'h9E},
{8'hFB, 8'hF3, 8'hC0},
{8'hF3, 8'hF1, 8'hC0},
{8'hF2, 8'hF3, 8'hDF},
{8'hF2, 8'hF2, 8'hE5},
{8'hE5, 8'hE5, 8'hDF},
{8'hDA, 8'hD8, 8'hD8},
{8'h85, 8'h83, 8'h87},
{8'h7E, 8'h7C, 8'h81},
{8'h7F, 8'h7D, 8'h81},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'h7F, 8'h7D, 8'h7E},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'h7C, 8'h7A, 8'h7D},
{8'h9B, 8'h9F, 8'h9B},
{8'hE9, 8'hF6, 8'hC8},
{8'hE7, 8'hF9, 8'hB5},
{8'hE1, 8'hF0, 8'hBE},
{8'hE1, 8'hF1, 8'hC3},
{8'hE1, 8'hF6, 8'hB4},
{8'hE1, 8'hF7, 8'hB2},
{8'hE1, 8'hF5, 8'hBF},
{8'hDD, 8'hEF, 8'hB3},
{8'hDF, 8'hEC, 8'hBC},
{8'hE4, 8'hE9, 8'hCE},
{8'hF2, 8'hF0, 8'hE8},
{8'hEE, 8'hE9, 8'hEB},
{8'hEF, 8'hEC, 8'hEE},
{8'hF2, 8'hF2, 8'hEC},
{8'hF3, 8'hF7, 8'hEC},
{8'hEA, 8'hEF, 8'hF6},
{8'hE8, 8'hEB, 8'hEC},
{8'hEF, 8'hEE, 8'hE5},
{8'hF8, 8'hF4, 8'hE9},
{8'hFD, 8'hF6, 8'hF5},
{8'hF9, 8'hF1, 8'hFD},
{8'hFA, 8'hF3, 8'hFF},
{8'hFE, 8'hFB, 8'hFF},
{8'hF9, 8'hF8, 8'hEB},
{8'hFB, 8'hF9, 8'hF1},
{8'hF5, 8'hF5, 8'hE7},
{8'hFA, 8'hF6, 8'hFA},
{8'hDE, 8'hD0, 8'hE6},
{8'hAC, 8'h9F, 8'h85},
{8'hE3, 8'hDB, 8'h9A},
{8'hBF, 8'hAA, 8'h8A},
{8'hEB, 8'hD2, 8'hBD},
{8'hAA, 8'h78, 8'h56},
{8'hF4, 8'hF7, 8'hB4},
{8'hFC, 8'hFC, 8'hB8},
{8'hCB, 8'h7B, 8'h5F},
{8'h76, 8'h34, 8'h34},
{8'h74, 8'h86, 8'h8B},
{8'h69, 8'h7B, 8'h8E},
{8'hB4, 8'hC1, 8'h9B},
{8'hFE, 8'hFF, 8'hCD},
{8'hC9, 8'hB8, 8'h99},
{8'h68, 8'h47, 8'h4E},
{8'hB9, 8'h98, 8'hA3},
{8'hFA, 8'hED, 8'hD4},
{8'hFF, 8'hFF, 8'hDA},
{8'hFB, 8'hFE, 8'hE0},
{8'hF1, 8'hFD, 8'hDF},
{8'hFF, 8'hFF, 8'hDE},
{8'hFF, 8'hE4, 8'hC7},
{8'hE4, 8'h8B, 8'h78},
{8'hB6, 8'h48, 8'h39},
{8'hAC, 8'h4B, 8'h34},
{8'hA9, 8'h61, 8'h38},
{8'hC7, 8'h93, 8'h58},
{8'h87, 8'h75, 8'h43},
{8'h29, 8'h42, 8'h76},
{8'h18, 8'h59, 8'hC5},
{8'h1F, 8'h55, 8'hAE},
{8'h24, 8'h2B, 8'h5C},
{8'h2F, 8'h1F, 8'h19},
{8'h28, 8'h21, 8'h17},
{8'h06, 8'h0D, 8'h2C},
{8'h00, 8'h18, 8'h24},
{8'h00, 8'h19, 8'h46},
{8'h06, 8'h12, 8'h6C},
{8'h09, 8'h17, 8'h7A},
{8'h25, 8'h31, 8'h75},
{8'h61, 8'h6E, 8'h83},
{8'hA1, 8'hAF, 8'hA0},
{8'hC1, 8'hCA, 8'hB0},
{8'hB7, 8'hBE, 8'hC0},
{8'hB8, 8'hBA, 8'hC0},
{8'hE8, 8'hE2, 8'hD5},
{8'hFD, 8'hF5, 8'hC8},
{8'hF9, 8'hEE, 8'hB4},
{8'hF9, 8'hEE, 8'hC0},
{8'hF8, 8'hF1, 8'hD3},
{8'hF8, 8'hF4, 8'hE0},
{8'hFA, 8'hFB, 8'hEB},
{8'hFA, 8'hFB, 8'hEE},
{8'hED, 8'hED, 8'hE7},
{8'h98, 8'h97, 8'h97},
{8'h7C, 8'h7A, 8'h7E},
{8'h7F, 8'h7D, 8'h82},
{8'hFF, 8'hD7, 8'h00},
{8'h7F, 8'h7D, 8'h7F},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'h7F, 8'h7C, 8'h83},
{8'h7F, 8'h7C, 8'h83},
{8'h7F, 8'h7D, 8'h82},
{8'h7F, 8'h7D, 8'h81},
{8'h7F, 8'h7D, 8'h82},
{8'h7F, 8'h7D, 8'h82},
{8'h7F, 8'h7C, 8'h82},
{8'h7C, 8'h79, 8'h81},
{8'hA8, 8'hAC, 8'hA6},
{8'hD6, 8'hE2, 8'hB3},
{8'hE8, 8'hF7, 8'hB6},
{8'hE1, 8'hEF, 8'hBE},
{8'hE3, 8'hF2, 8'hC5},
{8'hE2, 8'hF5, 8'hB4},
{8'hE1, 8'hF7, 8'hB0},
{8'hE2, 8'hF4, 8'hBE},
{8'hE2, 8'hF2, 8'hBF},
{8'hE2, 8'hED, 8'hC6},
{8'hD8, 8'hDB, 8'hC7},
{8'hF1, 8'hED, 8'hEA},
{8'hF8, 8'hF1, 8'hF6},
{8'hF7, 8'hF1, 8'hF7},
{8'hF5, 8'hF3, 8'hF2},
{8'hF3, 8'hF5, 8'hEF},
{8'hF1, 8'hF5, 8'hEF},
{8'hF5, 8'hF6, 8'hEF},
{8'hF6, 8'hF5, 8'hE6},
{8'hF9, 8'hF4, 8'hE1},
{8'hFC, 8'hF5, 8'hE2},
{8'hF9, 8'hF2, 8'hE7},
{8'hFB, 8'hF6, 8'hF2},
{8'hF9, 8'hF6, 8'hF3},
{8'hF4, 8'hF7, 8'hE7},
{8'hFA, 8'hFB, 8'hF2},
{8'hFA, 8'hF9, 8'hE1},
{8'hE6, 8'hE0, 8'hCE},
{8'h93, 8'h85, 8'h88},
{8'hA0, 8'h95, 8'h73},
{8'hE1, 8'hDA, 8'h99},
{8'hE7, 8'hDE, 8'hBC},
{8'hFF, 8'hFF, 8'hF6},
{8'hA5, 8'h9E, 8'h87},
{8'hB1, 8'hA7, 8'h7F},
{8'hFF, 8'hF9, 8'hC9},
{8'hFF, 8'hE9, 8'hBF},
{8'h9E, 8'h78, 8'h5B},
{8'h72, 8'h5F, 8'h50},
{8'h9B, 8'h8F, 8'h89},
{8'hEA, 8'hF5, 8'hBE},
{8'hF5, 8'hFD, 8'hC5},
{8'hA0, 8'h98, 8'h81},
{8'h18, 8'h04, 8'h0F},
{8'h20, 8'h00, 8'h12},
{8'h5A, 8'h3B, 8'h31},
{8'hC3, 8'hAA, 8'h86},
{8'hFC, 8'hF7, 8'hCF},
{8'hFF, 8'hFF, 8'hE1},
{8'hF2, 8'hD5, 8'hBB},
{8'hC8, 8'h70, 8'h64},
{8'hAA, 8'h30, 8'h27},
{8'h95, 8'h29, 8'h17},
{8'h8A, 8'h38, 8'h18},
{8'h9D, 8'h5C, 8'h32},
{8'hAE, 8'h76, 8'h47},
{8'h33, 8'h41, 8'h33},
{8'h12, 8'h51, 8'h9A},
{8'h13, 8'h54, 8'hB5},
{8'h16, 8'h22, 8'h59},
{8'h07, 8'h00, 8'h26},
{8'h00, 8'h02, 8'h34},
{8'h01, 8'h15, 8'h4C},
{8'h1B, 8'h1E, 8'h5D},
{8'h19, 8'h3A, 8'h80},
{8'h17, 8'h3E, 8'h9A},
{8'h1C, 8'h39, 8'hAE},
{8'h1B, 8'h36, 8'hAF},
{8'h19, 8'h31, 8'h98},
{8'h15, 8'h2E, 8'h7D},
{8'h1A, 8'h36, 8'h73},
{8'h45, 8'h5D, 8'h92},
{8'h99, 8'hA2, 8'hB4},
{8'hF8, 8'hFD, 8'hEC},
{8'hF8, 8'hFA, 8'hD1},
{8'hF6, 8'hF0, 8'hD1},
{8'hFE, 8'hF5, 8'hE3},
{8'hFE, 8'hF5, 8'hE3},
{8'hFA, 8'hF5, 8'hE9},
{8'hF6, 8'hF3, 8'hF4},
{8'hD8, 8'hD8, 8'hCD},
{8'hC4, 8'hC4, 8'hBB},
{8'h8C, 8'h8B, 8'h88},
{8'h7A, 8'h78, 8'h7B},
{8'h7F, 8'h7D, 8'h82},
{8'h7F, 8'h7D, 8'h82},
{8'hFF, 8'hD7, 8'h00},
{8'h7F, 8'h7D, 8'h7E},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'h7F, 8'h7C, 8'h85},
{8'h80, 8'h7D, 8'h85},
{8'h7F, 8'h7D, 8'h82},
{8'h82, 8'h80, 8'h82},
{8'h7F, 8'h7D, 8'h7F},
{8'h7F, 8'h7D, 8'h82},
{8'h7D, 8'h7A, 8'h82},
{8'h7E, 8'h7B, 8'h86},
{8'h7A, 8'h7D, 8'h77},
{8'hBD, 8'hC6, 8'h98},
{8'hEC, 8'hF9, 8'hBB},
{8'hE4, 8'hEF, 8'hC4},
{8'hE3, 8'hF0, 8'hC9},
{8'hE2, 8'hF4, 8'hB6},
{8'hE2, 8'hF7, 8'hB1},
{8'hE1, 8'hF3, 8'hBC},
{8'hE3, 8'hF1, 8'hBE},
{8'hE9, 8'hF2, 8'hC8},
{8'hE4, 8'hE6, 8'hCC},
{8'hE2, 8'hDE, 8'hD2},
{8'hF5, 8'hEF, 8'hEB},
{8'hF5, 8'hF0, 8'hED},
{8'hF8, 8'hF6, 8'hEF},
{8'hF9, 8'hFA, 8'hED},
{8'hF4, 8'hF9, 8'hE0},
{8'hFD, 8'hFD, 8'hEE},
{8'hF4, 8'hEF, 8'hEA},
{8'hFA, 8'hF0, 8'hEB},
{8'hFF, 8'hF7, 8'hE9},
{8'hFE, 8'hFA, 8'hE2},
{8'hF8, 8'hF4, 8'hDB},
{8'hF8, 8'hF6, 8'hE0},
{8'hF8, 8'hF9, 8'hF4},
{8'hFE, 8'hFD, 8'hFF},
{8'hDE, 8'hDE, 8'hBD},
{8'hDC, 8'hD9, 8'hA4},
{8'hDA, 8'hD0, 8'hAE},
{8'hB1, 8'hA5, 8'h78},
{8'hF1, 8'hE7, 8'hB1},
{8'hF3, 8'hE9, 8'hD1},
{8'hDF, 8'hDD, 8'hC2},
{8'hCD, 8'hA1, 8'h8C},
{8'h9F, 8'h57, 8'h43},
{8'hE3, 8'hB1, 8'h8B},
{8'hEE, 8'hDE, 8'hA4},
{8'hF2, 8'hF2, 8'hB7},
{8'hAF, 8'hA1, 8'h74},
{8'hCA, 8'hA3, 8'h8C},
{8'hFB, 8'hF3, 8'hC8},
{8'hF2, 8'hF3, 8'hCA},
{8'hF1, 8'hFA, 8'hE1},
{8'h97, 8'hA2, 8'h98},
{8'h1B, 8'h19, 8'h17},
{8'h16, 8'h00, 8'h00},
{8'h51, 8'h1D, 8'h0E},
{8'h99, 8'h5B, 8'h48},
{8'hBF, 8'h85, 8'h71},
{8'h7A, 8'h39, 8'h29},
{8'h67, 8'h27, 8'h1A},
{8'h62, 8'h25, 8'h11},
{8'h5B, 8'h1E, 8'h04},
{8'h6D, 8'h2E, 8'h0C},
{8'hA1, 8'h5F, 8'h3E},
{8'h82, 8'h41, 8'h2E},
{8'h18, 8'h2B, 8'h63},
{8'h1E, 8'h55, 8'hAB},
{8'h03, 8'h20, 8'h65},
{8'h02, 8'h00, 8'h15},
{8'h08, 8'h0B, 8'h26},
{8'h08, 8'h38, 8'h83},
{8'h18, 8'h53, 8'hBD},
{8'h31, 8'h4C, 8'hBA},
{8'h1F, 8'h50, 8'hC8},
{8'h1B, 8'h50, 8'hC2},
{8'h1E, 8'h54, 8'hBA},
{8'h1E, 8'h55, 8'hB1},
{8'h1A, 8'h52, 8'hAB},
{8'h1F, 8'h55, 8'hB5},
{8'h1A, 8'h4F, 8'hBE},
{8'h14, 8'h43, 8'hBA},
{8'h34, 8'h39, 8'h6B},
{8'hE3, 8'hEA, 8'hD8},
{8'hFE, 8'hFF, 8'hD6},
{8'hF4, 8'hF1, 8'hE2},
{8'hF7, 8'hF0, 8'hF6},
{8'hFB, 8'hF8, 8'hEF},
{8'hFC, 8'hFC, 8'hED},
{8'hF1, 8'hF1, 8'hF0},
{8'h89, 8'h89, 8'h81},
{8'h76, 8'h76, 8'h71},
{8'h7C, 8'h7A, 8'h7A},
{8'h84, 8'h82, 8'h86},
{8'h7F, 8'h7D, 8'h83},
{8'h7F, 8'h7D, 8'h82},
{8'h7F, 8'h7D, 8'h7F},
{8'h7F, 8'h7D, 8'h7D},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'h7F, 8'h7D, 8'h81},
{8'h7E, 8'h7B, 8'h86},
{8'h7E, 8'h7B, 8'h83},
{8'h80, 8'h7E, 8'h80},
{8'h81, 8'h80, 8'h7D},
{8'h7C, 8'h7B, 8'h78},
{8'h7E, 8'h7C, 8'h7E},
{8'h81, 8'h7E, 8'h85},
{8'h7F, 8'h7C, 8'h87},
{8'h97, 8'h99, 8'h95},
{8'hE7, 8'hEE, 8'hC5},
{8'hE6, 8'hF1, 8'hB9},
{8'hE3, 8'hEC, 8'hC9},
{8'hE2, 8'hEC, 8'hCC},
{8'hDC, 8'hEB, 8'hB4},
{8'hE4, 8'hF6, 8'hB5},
{8'hE6, 8'hF6, 8'hC1},
{8'hDF, 8'hED, 8'hB5},
{8'hE4, 8'hED, 8'hBC},
{8'hF0, 8'hF2, 8'hCE},
{8'hF3, 8'hF1, 8'hD9},
{8'hE3, 8'hDD, 8'hCD},
{8'hEA, 8'hE5, 8'hD5},
{8'hE3, 8'hE1, 8'hCF},
{8'hF6, 8'hF8, 8'hE3},
{8'hF9, 8'hF7, 8'hF5},
{8'hF0, 8'hEB, 8'hF1},
{8'hF1, 8'hE7, 8'hED},
{8'hF9, 8'hEE, 8'hE4},
{8'hF7, 8'hEE, 8'hCF},
{8'hF9, 8'hF2, 8'hCE},
{8'hF9, 8'hF2, 8'hDF},
{8'hFA, 8'hF3, 8'hF1},
{8'hF4, 8'hF6, 8'hEC},
{8'hBC, 8'hBD, 8'hCB},
{8'hAB, 8'hAD, 8'hA5},
{8'hB6, 8'hBA, 8'h9A},
{8'hBB, 8'hB8, 8'hAA},
{8'hB4, 8'hA6, 8'h90},
{8'hD1, 8'hC2, 8'h91},
{8'h8D, 8'h75, 8'h51},
{8'h85, 8'h50, 8'h1F},
{8'hBE, 8'h46, 8'h2C},
{8'hA7, 8'h4A, 8'h34},
{8'h98, 8'h68, 8'h40},
{8'hDD, 8'hAA, 8'h79},
{8'hC0, 8'hB5, 8'h73},
{8'hE0, 8'hF2, 8'hB9},
{8'hEC, 8'hD3, 8'hB7},
{8'hF2, 8'hEB, 8'hD2},
{8'hF7, 8'hF8, 8'hE5},
{8'hF4, 8'hFC, 8'hE9},
{8'hEF, 8'hFA, 8'hE0},
{8'hD4, 8'hD7, 8'hC1},
{8'h78, 8'h61, 8'h5C},
{8'h49, 8'h15, 8'h1A},
{8'h5E, 8'h16, 8'h17},
{8'h6C, 8'h0D, 8'h07},
{8'h4B, 8'h16, 8'h0F},
{8'h26, 8'h1C, 8'h11},
{8'h1F, 8'h1A, 8'h09},
{8'h36, 8'h17, 8'h02},
{8'h67, 8'h31, 8'h15},
{8'h92, 8'h5E, 8'h4A},
{8'h3B, 8'h1D, 8'h1D},
{8'h16, 8'h32, 8'h85},
{8'h10, 8'h22, 8'h64},
{8'h01, 8'h00, 8'h2F},
{8'h03, 8'h08, 8'h36},
{8'h16, 8'h3D, 8'h75},
{8'h16, 8'h5C, 8'hB4},
{8'h08, 8'h52, 8'hC1},
{8'h16, 8'h58, 8'hC1},
{8'h13, 8'h59, 8'hAE},
{8'h10, 8'h58, 8'hA7},
{8'h0F, 8'h58, 8'hA3},
{8'h0F, 8'h5A, 8'hA8},
{8'h0F, 8'h59, 8'hB0},
{8'h0C, 8'h57, 8'hB3},
{8'h0A, 8'h57, 8'hB1},
{8'h0F, 8'h57, 8'hAD},
{8'h24, 8'h26, 8'h5D},
{8'hDE, 8'hE0, 8'hDE},
{8'hFA, 8'hFD, 8'hE2},
{8'hF9, 8'hF8, 8'hF2},
{8'hF5, 8'hF2, 8'hF8},
{8'hF0, 8'hF0, 8'hE3},
{8'hFD, 8'hFE, 8'hE5},
{8'hF1, 8'hF3, 8'hE3},
{8'hA3, 8'hA3, 8'h9D},
{8'h7F, 8'h7E, 8'h7B},
{8'h81, 8'h7F, 8'h82},
{8'h7B, 8'h79, 8'h7F},
{8'h7E, 8'h7B, 8'h82},
{8'h7F, 8'h7D, 8'h82},
{8'h7F, 8'h7D, 8'h7F},
{8'h7F, 8'h7E, 8'h7C},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'h80, 8'h7E, 8'h81},
{8'h82, 8'h7F, 8'h88},
{8'h79, 8'h77, 8'h7B},
{8'h7D, 8'h7C, 8'h77},
{8'h82, 8'h82, 8'h77},
{8'h85, 8'h84, 8'h7A},
{8'h79, 8'h78, 8'h74},
{8'hFF, 8'hD7, 8'h00},
{8'h78, 8'h75, 8'h7F},
{8'h9C, 8'h9B, 8'h9C},
{8'hEA, 8'hF0, 8'hCC},
{8'hE9, 8'hF2, 8'hC3},
{8'hB5, 8'hBA, 8'hA1},
{8'h89, 8'h91, 8'h7D},
{8'hCE, 8'hDA, 8'hAC},
{8'hE6, 8'hF5, 8'hBA},
{8'hE2, 8'hF0, 8'hC0},
{8'hE1, 8'hED, 8'hB9},
{8'hE6, 8'hED, 8'hBE},
{8'hF2, 8'hF4, 8'hCE},
{8'hFD, 8'hFA, 8'hDF},
{8'hE7, 8'hE1, 8'hCC},
{8'hE9, 8'hE3, 8'hD0},
{8'hD8, 8'hD6, 8'hC1},
{8'hED, 8'hEC, 8'hD8},
{8'hF4, 8'hF0, 8'hF0},
{8'hF3, 8'hEC, 8'hE8},
{8'hF2, 8'hEA, 8'hCC},
{8'hF0, 8'hEC, 8'hA3},
{8'hE5, 8'hE4, 8'h7C},
{8'hE9, 8'hE9, 8'h8A},
{8'hF5, 8'hEF, 8'hC2},
{8'hF9, 8'hF1, 8'hEC},
{8'hBC, 8'hCB, 8'hBC},
{8'h2F, 8'h3E, 8'h66},
{8'h13, 8'h27, 8'h57},
{8'h04, 8'h18, 8'h3A},
{8'h01, 8'h09, 8'h39},
{8'h31, 8'h2C, 8'h45},
{8'h85, 8'h78, 8'h56},
{8'hC4, 8'hA8, 8'h6F},
{8'hDD, 8'hA7, 8'h8D},
{8'h76, 8'h3C, 8'h38},
{8'h2B, 8'h0E, 8'h10},
{8'h4F, 8'h32, 8'h26},
{8'hAF, 8'h6C, 8'h4B},
{8'hC4, 8'h83, 8'h48},
{8'hB1, 8'h90, 8'h4A},
{8'hF2, 8'hE1, 8'hA6},
{8'hC3, 8'hCA, 8'hAE},
{8'hCC, 8'hD0, 8'hCB},
{8'hFE, 8'hFD, 8'hF9},
{8'hFF, 8'hFD, 8'hE8},
{8'hFF, 8'hFF, 8'hF3},
{8'hCD, 8'hB5, 8'hBE},
{8'h29, 8'h08, 8'h12},
{8'h3B, 8'h14, 8'h0F},
{8'h49, 8'h11, 8'h09},
{8'h18, 8'h02, 8'h04},
{8'h00, 8'h02, 8'h0A},
{8'h00, 8'h01, 8'h03},
{8'h34, 8'h18, 8'h10},
{8'h57, 8'h2B, 8'h21},
{8'h5D, 8'h45, 8'h3F},
{8'h07, 8'h0A, 8'h16},
{8'h1C, 8'h2F, 8'h6E},
{8'h04, 8'h02, 8'h1C},
{8'h07, 8'h00, 8'h2B},
{8'h12, 8'h2A, 8'h83},
{8'h19, 8'h57, 8'hB6},
{8'h16, 8'h5A, 8'hBB},
{8'h13, 8'h58, 8'hB7},
{8'h08, 8'h57, 8'hA2},
{8'h12, 8'h55, 8'hB8},
{8'h14, 8'h59, 8'hB3},
{8'h13, 8'h5A, 8'hAB},
{8'h0F, 8'h56, 8'hAD},
{8'h10, 8'h56, 8'hBD},
{8'h0D, 8'h52, 8'hC0},
{8'h0F, 8'h58, 8'hBF},
{8'h0C, 8'h50, 8'hA9},
{8'h1D, 8'h1C, 8'h3D},
{8'hEC, 8'hE8, 8'hEE},
{8'hFE, 8'hFD, 8'hFB},
{8'hFB, 8'hFA, 8'hF5},
{8'hF3, 8'hF3, 8'hEA},
{8'hDD, 8'hDF, 8'hCB},
{8'hD9, 8'hDC, 8'hC0},
{8'hAF, 8'hB2, 8'h99},
{8'h7A, 8'h78, 8'h75},
{8'h7D, 8'h7C, 8'h7D},
{8'h7D, 8'h7A, 8'h80},
{8'h81, 8'h7E, 8'h86},
{8'h7F, 8'h7C, 8'h84},
{8'h7F, 8'h7D, 8'h81},
{8'h7F, 8'h7E, 8'h7E},
{8'h7F, 8'h7E, 8'h7B},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'h81, 8'h7E, 8'h85},
{8'h7C, 8'h7B, 8'h7B},
{8'h7A, 8'h7A, 8'h6F},
{8'h96, 8'h97, 8'h85},
{8'hD3, 8'hD4, 8'hC3},
{8'h91, 8'h90, 8'h87},
{8'h76, 8'h75, 8'h75},
{8'h7B, 8'h77, 8'h80},
{8'h7D, 8'h7A, 8'h80},
{8'hB0, 8'hB4, 8'h96},
{8'hEC, 8'hF2, 8'hCA},
{8'h97, 8'h9B, 8'h8B},
{8'h80, 8'h84, 8'h79},
{8'hD9, 8'hE4, 8'hBD},
{8'hE4, 8'hF1, 8'hBC},
{8'hE4, 8'hF1, 8'hC6},
{8'hE2, 8'hEB, 8'hC3},
{8'hDE, 8'hE3, 8'hBF},
{8'hEB, 8'hEA, 8'hCE},
{8'hFD, 8'hFB, 8'hE8},
{8'hF4, 8'hED, 8'hDF},
{8'hD8, 8'hD0, 8'hC4},
{8'hF3, 8'hEE, 8'hE2},
{8'hF5, 8'hF3, 8'hE6},
{8'hF2, 8'hEE, 8'hE1},
{8'hF9, 8'hF3, 8'hE5},
{8'hF4, 8'hEC, 8'hCA},
{8'hE6, 8'hE1, 8'h92},
{8'hDC, 8'hDD, 8'h66},
{8'hD4, 8'hD6, 8'h62},
{8'hEF, 8'hEA, 8'hA9},
{8'hFD, 8'hF7, 8'hE6},
{8'h5A, 8'h78, 8'h8B},
{8'h22, 8'h48, 8'hA1},
{8'h1C, 8'h54, 8'hB5},
{8'h1A, 8'h5C, 8'hA5},
{8'h15, 8'h46, 8'h9B},
{8'h14, 8'h23, 8'h64},
{8'h33, 8'h28, 8'h28},
{8'h5E, 8'h41, 8'h27},
{8'h2B, 8'h1F, 8'h23},
{8'h10, 8'h1D, 8'h39},
{8'h08, 8'h1E, 8'h4A},
{8'h24, 8'h22, 8'h40},
{8'h56, 8'h26, 8'h20},
{8'hAD, 8'h5F, 8'h3D},
{8'h94, 8'h51, 8'h24},
{8'hC4, 8'h97, 8'h68},
{8'hE0, 8'hDC, 8'hB4},
{8'h49, 8'h45, 8'h44},
{8'h95, 8'h93, 8'h9F},
{8'hB4, 8'hB8, 8'hB5},
{8'h94, 8'h96, 8'h97},
{8'h53, 8'h47, 8'h5D},
{8'h16, 8'h02, 8'h07},
{8'h3C, 8'h1E, 8'h05},
{8'h26, 8'h19, 8'h0D},
{8'h07, 8'h00, 8'h0E},
{8'h06, 8'h00, 8'h22},
{8'h06, 8'h00, 8'h15},
{8'h29, 8'h1C, 8'h1A},
{8'h3B, 8'h2B, 8'h26},
{8'h26, 8'h1D, 8'h27},
{8'h10, 8'h0B, 8'h33},
{8'h0F, 8'h12, 8'h44},
{8'h04, 8'h02, 8'h0E},
{8'h05, 8'h0C, 8'h32},
{8'h1C, 8'h4A, 8'h9F},
{8'h11, 8'h5A, 8'hB0},
{8'h16, 8'h56, 8'hB5},
{8'h20, 8'h50, 8'hB3},
{8'h1D, 8'h51, 8'h94},
{8'h1C, 8'h4E, 8'hB9},
{8'h18, 8'h4D, 8'hAA},
{8'h18, 8'h50, 8'h9F},
{8'h1D, 8'h54, 8'hAC},
{8'h1B, 8'h4F, 8'hBA},
{8'h1B, 8'h4F, 8'hC1},
{8'h1E, 8'h54, 8'hBA},
{8'h01, 8'h30, 8'h81},
{8'h37, 8'h34, 8'h34},
{8'hF8, 8'hF1, 8'hF5},
{8'hFF, 8'hFC, 8'hFF},
{8'hE8, 8'hE8, 8'hDC},
{8'hD5, 8'hD8, 8'hBB},
{8'hA9, 8'hAA, 8'h97},
{8'h75, 8'h73, 8'h68},
{8'h84, 8'h83, 8'h74},
{8'h79, 8'h77, 8'h78},
{8'h7D, 8'h7B, 8'h80},
{8'h81, 8'h7E, 8'h85},
{8'h7E, 8'h7A, 8'h84},
{8'h7F, 8'h7B, 8'h84},
{8'h7F, 8'h7D, 8'h81},
{8'h7F, 8'h7E, 8'h7D},
{8'h7F, 8'h7E, 8'h7A},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'h7F, 8'h7E, 8'h7F},
{8'h85, 8'h86, 8'h7E},
{8'h7E, 8'h7E, 8'h78},
{8'h7F, 8'h80, 8'h7A},
{8'h7D, 8'h7E, 8'h72},
{8'hC2, 8'hC5, 8'hB3},
{8'hE0, 8'hE3, 8'hD1},
{8'h8D, 8'h90, 8'h84},
{8'h7C, 8'h7D, 8'h7B},
{8'h7D, 8'h7C, 8'h83},
{8'h7E, 8'h81, 8'h6C},
{8'h95, 8'h9A, 8'h7C},
{8'h7A, 8'h7C, 8'h6F},
{8'hC0, 8'hC3, 8'hB8},
{8'hAF, 8'hB7, 8'h97},
{8'hD0, 8'hD9, 8'hAF},
{8'hE5, 8'hED, 8'hCB},
{8'hE8, 8'hEC, 8'hD2},
{8'hF1, 8'hF3, 8'hDC},
{8'hF7, 8'hF5, 8'hE3},
{8'hF5, 8'hEE, 8'hE3},
{8'hEB, 8'hE4, 8'hDD},
{8'hF0, 8'hE9, 8'hE6},
{8'hFD, 8'hF8, 8'hF5},
{8'hF9, 8'hF6, 8'hF4},
{8'hFA, 8'hF4, 8'hF2},
{8'hFA, 8'hF0, 8'hF7},
{8'hFD, 8'hF0, 8'hF2},
{8'hFF, 8'hF6, 8'hDD},
{8'hF4, 8'hEB, 8'hAF},
{8'hE8, 8'hE0, 8'h9C},
{8'hF8, 8'hEE, 8'hC4},
{8'hDC, 8'hD1, 8'hC7},
{8'h1F, 8'h3B, 8'h75},
{8'h24, 8'h55, 8'hC5},
{8'h0E, 8'h52, 8'hBD},
{8'h0C, 8'h5D, 8'hA9},
{8'h18, 8'h5C, 8'hB3},
{8'h23, 8'h4A, 8'h9C},
{8'h19, 8'h20, 8'h4C},
{8'h30, 8'h2A, 8'h3E},
{8'h04, 8'h16, 8'h19},
{8'h03, 8'h02, 8'h21},
{8'h06, 8'h1D, 8'h4D},
{8'h23, 8'h39, 8'h68},
{8'h21, 8'h06, 8'h1E},
{8'h5E, 8'h3A, 8'h34},
{8'h27, 8'h15, 8'h0C},
{8'h60, 8'h2F, 8'h30},
{8'hE2, 8'hBE, 8'h9B},
{8'h8B, 8'h7A, 8'h7E},
{8'h18, 8'h25, 8'h44},
{8'h03, 8'h1A, 8'h34},
{8'h00, 8'h00, 8'h1B},
{8'h00, 8'h00, 8'h19},
{8'h22, 8'h06, 8'h0A},
{8'h45, 8'h21, 8'h00},
{8'h12, 8'h17, 8'h08},
{8'h04, 8'h00, 8'h0C},
{8'h09, 8'h01, 8'h27},
{8'h05, 8'h10, 8'h38},
{8'h17, 8'h2D, 8'h48},
{8'h15, 8'h20, 8'h2F},
{8'h09, 8'h02, 8'h1E},
{8'h19, 8'h01, 8'h35},
{8'h07, 8'h01, 8'h2C},
{8'h00, 8'h01, 8'h14},
{8'h0C, 8'h23, 8'h4C},
{8'h21, 8'h59, 8'h9D},
{8'h11, 8'h58, 8'h97},
{8'h04, 8'h34, 8'h88},
{8'h11, 8'h2E, 8'h96},
{8'h24, 8'h42, 8'h93},
{8'h13, 8'h4B, 8'h8F},
{8'h08, 8'h35, 8'h77},
{8'h0E, 8'h28, 8'h65},
{8'h0E, 8'h21, 8'h67},
{8'h18, 8'h34, 8'h89},
{8'h2E, 8'h4D, 8'hA2},
{8'h24, 8'h4B, 8'h80},
{8'h12, 8'h33, 8'h41},
{8'h7C, 8'h7B, 8'h65},
{8'hE4, 8'hD9, 8'hD7},
{8'hED, 8'hDB, 8'hE6},
{8'hF8, 8'hF0, 8'hE5},
{8'hD1, 8'hD3, 8'hB1},
{8'h7E, 8'h80, 8'h6C},
{8'hBD, 8'hBC, 8'hB3},
{8'hED, 8'hEA, 8'hDC},
{8'hCF, 8'hCC, 8'hC5},
{8'h96, 8'h97, 8'h95},
{8'h78, 8'h7C, 8'h80},
{8'h7B, 8'h7F, 8'h85},
{8'h7B, 8'h7C, 8'h82},
{8'h80, 8'h7D, 8'h81},
{8'h81, 8'h7C, 8'h7F},
{8'h81, 8'h7C, 8'h7F},
{8'h7F, 8'h7D, 8'h7E},
{8'h7F, 8'h7D, 8'h7E},
{8'h80, 8'h7E, 8'h80},
{8'h7F, 8'h7D, 8'h7F},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'h80, 8'h7F, 8'h7D},
{8'hC3, 8'hCB, 8'h9F},
{8'hB0, 8'hB4, 8'hA3},
{8'h75, 8'h76, 8'h82},
{8'h76, 8'h79, 8'h85},
{8'h8A, 8'h92, 8'h84},
{8'hE4, 8'hF1, 8'hCB},
{8'hD8, 8'hE7, 8'hBD},
{8'h93, 8'hA0, 8'h7F},
{8'h76, 8'h7A, 8'h7A},
{8'h77, 8'h7A, 8'h78},
{8'h76, 8'h79, 8'h6F},
{8'h91, 8'h95, 8'h83},
{8'hD4, 8'hD6, 8'hC1},
{8'hB9, 8'hBA, 8'hA7},
{8'hE0, 8'hE0, 8'hD1},
{8'hF6, 8'hF4, 8'hE8},
{8'hF1, 8'hED, 8'hE0},
{8'hF8, 8'hF4, 8'hE7},
{8'hF2, 8'hEF, 8'hE1},
{8'hE0, 8'hDF, 8'hD3},
{8'hED, 8'hEC, 8'hE5},
{8'hF7, 8'hF8, 8'hF8},
{8'hF9, 8'hF8, 8'hFD},
{8'hF3, 8'hF2, 8'hFD},
{8'hF6, 8'hF5, 8'hF8},
{8'hF4, 8'hF5, 8'hEE},
{8'hFA, 8'hFA, 8'hE8},
{8'hEE, 8'hED, 8'hCF},
{8'hEC, 8'hE9, 8'hC8},
{8'hF2, 8'hEB, 8'hCD},
{8'hFF, 8'hFB, 8'hE3},
{8'h96, 8'h91, 8'h87},
{8'h0F, 8'h3A, 8'h82},
{8'h1E, 8'h53, 8'hA3},
{8'h1A, 8'h51, 8'hA4},
{8'h1C, 8'h56, 8'hAD},
{8'h18, 8'h56, 8'hAD},
{8'h1C, 8'h59, 8'hAF},
{8'h15, 8'h4E, 8'hA4},
{8'h10, 8'h46, 8'h9A},
{8'h25, 8'h43, 8'h7D},
{8'h03, 8'h0F, 8'h33},
{8'h02, 8'h06, 8'h30},
{8'h38, 8'h34, 8'h76},
{8'h0B, 8'h06, 8'h37},
{8'h1E, 8'h1D, 8'h22},
{8'h14, 8'h17, 8'h0D},
{8'h00, 8'h00, 8'h03},
{8'h71, 8'h51, 8'h5E},
{8'h92, 8'h9E, 8'h9F},
{8'h20, 8'h56, 8'h8D},
{8'h1E, 8'h4F, 8'hCB},
{8'h25, 8'h39, 8'h87},
{8'h4B, 8'h4D, 8'h31},
{8'h31, 8'h26, 8'h09},
{8'h19, 8'h0E, 8'h38},
{8'h08, 8'h1D, 8'h39},
{8'h10, 8'h27, 8'h46},
{8'h18, 8'h3B, 8'h7B},
{8'h0F, 8'h50, 8'hB7},
{8'h12, 8'h48, 8'hB0},
{8'h02, 8'h09, 8'h46},
{8'h0A, 8'h00, 8'h1B},
{8'h09, 8'h01, 8'h12},
{8'h06, 8'h03, 8'h0A},
{8'h00, 8'h01, 8'h2A},
{8'h14, 8'h2A, 8'h79},
{8'h22, 8'h52, 8'hAF},
{8'h0E, 8'h47, 8'h9A},
{8'h13, 8'h4A, 8'h92},
{8'h22, 8'h55, 8'hA4},
{8'h1F, 8'h48, 8'hA2},
{8'h03, 8'h42, 8'h90},
{8'h08, 8'h46, 8'h99},
{8'h14, 8'h42, 8'h8F},
{8'h16, 8'h33, 8'h71},
{8'h0D, 8'h17, 8'h4F},
{8'h1C, 8'h20, 8'h53},
{8'h7D, 8'h88, 8'h9C},
{8'hD0, 8'hDF, 8'hD2},
{8'hFC, 8'hFF, 8'hE6},
{8'hFD, 8'hF7, 8'hE6},
{8'hFA, 8'hE5, 8'hDD},
{8'hEB, 8'hD6, 8'hCC},
{8'hE4, 8'hE7, 8'hD2},
{8'hB7, 8'hC8, 8'hA7},
{8'hDB, 8'hE3, 8'hBD},
{8'hE5, 8'hDE, 8'hB7},
{8'hE7, 8'hD5, 8'hB2},
{8'hB3, 8'hB2, 8'h9B},
{8'h70, 8'h82, 8'h77},
{8'h6F, 8'h84, 8'h80},
{8'h79, 8'h83, 8'h7F},
{8'h7B, 8'h76, 8'h77},
{8'h84, 8'h76, 8'h82},
{8'h85, 8'h76, 8'h8A},
{8'h7C, 8'h7B, 8'h78},
{8'h85, 8'h84, 8'h80},
{8'h82, 8'h81, 8'h7F},
{8'h7E, 8'h7D, 8'h7C},
{8'h7F, 8'h7D, 8'h7F},
{8'hFF, 8'hD7, 8'h00},
{8'h7F, 8'h7D, 8'h81},
{8'h7F, 8'h7D, 8'h82},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'h7B, 8'h79, 8'h7A},
{8'hA4, 8'hA9, 8'h8F},
{8'hEB, 8'hF0, 8'hDB},
{8'hAE, 8'hB2, 8'hA6},
{8'h79, 8'h80, 8'h72},
{8'h75, 8'h7E, 8'h66},
{8'hC1, 8'hCF, 8'hAA},
{8'hE6, 8'hF4, 8'hC9},
{8'hD8, 8'hE7, 8'hBD},
{8'h9E, 8'hA4, 8'h9B},
{8'h76, 8'h7B, 8'h71},
{8'h87, 8'h8B, 8'h7C},
{8'hD7, 8'hDB, 8'hC9},
{8'hC8, 8'hCA, 8'hB7},
{8'hCA, 8'hCB, 8'hBB},
{8'hFF, 8'hFF, 8'hF5},
{8'hF5, 8'hF2, 8'hEC},
{8'hF2, 8'hED, 8'hE6},
{8'hE4, 8'hE0, 8'hD7},
{8'hD5, 8'hD2, 8'hC6},
{8'hE8, 8'hE7, 8'hDA},
{8'hFA, 8'hFA, 8'hED},
{8'hF9, 8'hFA, 8'hF2},
{8'hFB, 8'hFB, 8'hF8},
{8'hFA, 8'hFB, 8'hF9},
{8'hF5, 8'hFC, 8'hF3},
{8'hF1, 8'hF7, 8'hE9},
{8'hEF, 8'hF6, 8'hDE},
{8'hE1, 8'hE9, 8'hCA},
{8'hEF, 8'hF4, 8'hD5},
{8'hF6, 8'hFB, 8'hE1},
{8'hF4, 8'hF7, 8'hE4},
{8'h52, 8'h56, 8'h56},
{8'h02, 8'h40, 8'h9B},
{8'h0E, 8'h58, 8'hB9},
{8'h12, 8'h5A, 8'hBA},
{8'h13, 8'h58, 8'hB5},
{8'h1E, 8'h5D, 8'hB6},
{8'h1A, 8'h51, 8'hA4},
{8'h25, 8'h56, 8'hA1},
{8'h27, 8'h53, 8'h9F},
{8'h20, 8'h56, 8'hB9},
{8'h16, 8'h41, 8'h8E},
{8'h00, 8'h0C, 8'h47},
{8'h21, 8'h22, 8'h5E},
{8'h1B, 8'h1A, 8'h54},
{8'h09, 8'h0F, 8'h3F},
{8'h09, 8'h23, 8'h45},
{8'h02, 8'h18, 8'h35},
{8'h0B, 8'h1E, 8'h49},
{8'h44, 8'h73, 8'h9D},
{8'h1B, 8'h53, 8'h9E},
{8'h34, 8'h59, 8'hAA},
{8'h69, 8'h78, 8'h68},
{8'hDF, 8'hE8, 8'h73},
{8'h89, 8'h8F, 8'h53},
{8'h35, 8'h39, 8'h87},
{8'h25, 8'h40, 8'hC2},
{8'h24, 8'h4C, 8'hC8},
{8'h12, 8'h54, 8'hCC},
{8'h0F, 8'h59, 8'hBD},
{8'h1E, 8'h42, 8'h75},
{8'h0F, 8'h05, 8'h09},
{8'h0B, 8'h00, 8'h01},
{8'h00, 8'h09, 8'h1E},
{8'h05, 8'h05, 8'h12},
{8'h01, 8'h06, 8'h2E},
{8'h1E, 8'h39, 8'h85},
{8'h1E, 8'h4F, 8'hA9},
{8'h19, 8'h57, 8'hAC},
{8'h18, 8'h57, 8'hA4},
{8'h18, 8'h49, 8'h9B},
{8'h08, 8'h21, 8'h7B},
{8'h13, 8'h24, 8'h70},
{8'h11, 8'h4F, 8'h92},
{8'h03, 8'h5C, 8'hB4},
{8'h09, 8'h56, 8'hC8},
{8'h2B, 8'h50, 8'hAA},
{8'h76, 8'h7A, 8'h97},
{8'hF6, 8'hF0, 8'hEE},
{8'hFF, 8'hFB, 8'hFF},
{8'hF7, 8'hFC, 8'hE3},
{8'hFA, 8'hF9, 8'hE2},
{8'hF5, 8'hF4, 8'hE0},
{8'hF2, 8'hF8, 8'hE4},
{8'hE2, 8'hF1, 8'hD7},
{8'hE7, 8'hF1, 8'hD1},
{8'hEB, 8'hE0, 8'hC3},
{8'hED, 8'hCC, 8'hB3},
{8'hEF, 8'hC0, 8'hA6},
{8'hB4, 8'h94, 8'h80},
{8'h7E, 8'h76, 8'h6A},
{8'h7B, 8'h7E, 8'h73},
{8'h90, 8'h93, 8'h83},
{8'h95, 8'h93, 8'h83},
{8'h84, 8'h82, 8'h78},
{8'h7C, 8'h7D, 8'h7A},
{8'h7F, 8'h7F, 8'h7B},
{8'h95, 8'h94, 8'h91},
{8'h7F, 8'h7E, 8'h7C},
{8'h7C, 8'h7A, 8'h7A},
{8'h7F, 8'h7D, 8'h7F},
{8'hFF, 8'hD7, 8'h00},
{8'h7F, 8'h7D, 8'h81},
{8'h7F, 8'h7D, 8'h82},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'h7C, 8'h7E, 8'h79},
{8'hCC, 8'hD1, 8'hBA},
{8'hEC, 8'hF6, 8'hCC},
{8'hAF, 8'hBA, 8'h8D},
{8'h82, 8'h8E, 8'h68},
{8'hC3, 8'hD0, 8'hAB},
{8'hE5, 8'hF5, 8'hC5},
{8'hDF, 8'hF1, 8'hB7},
{8'hE6, 8'hF0, 8'hD1},
{8'hBA, 8'hC2, 8'hA5},
{8'h9C, 8'hA2, 8'h85},
{8'hAC, 8'hB2, 8'h96},
{8'hD0, 8'hD3, 8'hBC},
{8'hDD, 8'hDE, 8'hCD},
{8'hCB, 8'hCA, 8'hBF},
{8'hE5, 8'hE2, 8'hDB},
{8'hF7, 8'hF2, 8'hF3},
{8'hED, 8'hE7, 8'hE5},
{8'hE1, 8'hDE, 8'hD6},
{8'hEA, 8'hE9, 8'hDB},
{8'hF2, 8'hF4, 8'hE0},
{8'hF1, 8'hF3, 8'hDF},
{8'hEB, 8'hEE, 8'hDB},
{8'hDF, 8'hE1, 8'hD1},
{8'hE7, 8'hD9, 8'hDA},
{8'hEC, 8'hDE, 8'hDC},
{8'hE8, 8'hDC, 8'hD7},
{8'hF9, 8'hF3, 8'hEC},
{8'hFA, 8'hF3, 8'hF2},
{8'hFA, 8'hF3, 8'hFA},
{8'hF2, 8'hEB, 8'hF2},
{8'h2A, 8'h29, 8'h43},
{8'h0E, 8'h4C, 8'hA4},
{8'h16, 8'h59, 8'hB5},
{8'h1B, 8'h5A, 8'hB2},
{8'h0F, 8'h43, 8'h95},
{8'h0A, 8'h2C, 8'h78},
{8'h05, 8'h15, 8'h57},
{8'h0A, 8'h14, 8'h4D},
{8'h10, 8'h22, 8'h56},
{8'h0C, 8'h37, 8'h7A},
{8'h21, 8'h4C, 8'h9E},
{8'h0D, 8'h2A, 8'h70},
{8'h0B, 8'h23, 8'h44},
{8'h13, 8'h32, 8'h4B},
{8'h01, 8'h11, 8'h4E},
{8'h21, 8'h3B, 8'hA3},
{8'h1F, 8'h34, 8'hA5},
{8'h1A, 8'h1E, 8'h49},
{8'h55, 8'h5F, 8'h6D},
{8'h8E, 8'h91, 8'h81},
{8'hC4, 8'hB1, 8'h83},
{8'hEC, 8'hBA, 8'h6B},
{8'hF0, 8'hBD, 8'h5A},
{8'hF0, 8'hD4, 8'h76},
{8'hC8, 8'hBD, 8'h77},
{8'h83, 8'h90, 8'h97},
{8'h56, 8'h69, 8'h81},
{8'h2A, 8'h55, 8'h8B},
{8'h1C, 8'h5B, 8'hA8},
{8'h14, 8'h3B, 8'h7A},
{8'h05, 8'h02, 8'h1D},
{8'h03, 8'h01, 8'h10},
{8'h00, 8'h0A, 8'h26},
{8'h05, 8'h05, 8'h17},
{8'h03, 8'h08, 8'h2F},
{8'h1C, 8'h39, 8'h7F},
{8'h1D, 8'h4D, 8'hA3},
{8'h17, 8'h53, 8'hAB},
{8'h17, 8'h55, 8'hA9},
{8'h06, 8'h2F, 8'h85},
{8'h12, 8'h3B, 8'h97},
{8'h2F, 8'h45, 8'hA9},
{8'h1B, 8'h55, 8'hB8},
{8'h07, 8'h5E, 8'hC1},
{8'h17, 8'h5D, 8'hB4},
{8'h51, 8'h68, 8'h94},
{8'hE0, 8'hD6, 8'hD2},
{8'hFF, 8'hF9, 8'hE6},
{8'hF9, 8'hF9, 8'hEE},
{8'hFD, 8'hF6, 8'hDF},
{8'hFF, 8'hF4, 8'hDA},
{8'hFD, 8'hF5, 8'hDC},
{8'hFA, 8'hF5, 8'hDA},
{8'hFB, 8'hF6, 8'hD8},
{8'hF7, 8'hD8, 8'hBD},
{8'hF6, 8'hB5, 8'hA0},
{8'hFA, 8'hA3, 8'h92},
{8'hE3, 8'h9B, 8'h80},
{8'hBD, 8'h8D, 8'h77},
{8'hBB, 8'hA6, 8'h92},
{8'hDC, 8'hD8, 8'hC0},
{8'hEF, 8'hF0, 8'hCC},
{8'hF1, 8'hF2, 8'hCB},
{8'hDB, 8'hE2, 8'hBF},
{8'h99, 8'hA7, 8'h8B},
{8'h8E, 8'h8F, 8'h89},
{8'h95, 8'h94, 8'h91},
{8'h7E, 8'h7D, 8'h7B},
{8'h7C, 8'h7A, 8'h7A},
{8'h7F, 8'h7D, 8'h7F},
{8'hFF, 8'hD7, 8'h00},
{8'h7F, 8'h7D, 8'h81},
{8'h7F, 8'h7D, 8'h82},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'h7E, 8'h7C, 8'h80},
{8'h78, 8'h78, 8'h81},
{8'hA1, 8'hA6, 8'h8F},
{8'hE8, 8'hF5, 8'hBA},
{8'hE8, 8'hF6, 8'hB6},
{8'hD8, 8'hE6, 8'hB5},
{8'hE0, 8'hEE, 8'hC7},
{8'hE4, 8'hF5, 8'hC0},
{8'hE3, 8'hF6, 8'hB2},
{8'hE3, 8'hF1, 8'hB8},
{8'hE4, 8'hF0, 8'hBA},
{8'hE7, 8'hEF, 8'hC0},
{8'hD8, 8'hE0, 8'hB5},
{8'hE1, 8'hE5, 8'hC3},
{8'hE5, 8'hE7, 8'hCC},
{8'hA0, 8'hA0, 8'h8B},
{8'hC0, 8'hBF, 8'hAE},
{8'hFD, 8'hF9, 8'hFD},
{8'hFD, 8'hF9, 8'hFA},
{8'hF6, 8'hF2, 8'hEC},
{8'hDE, 8'hDD, 8'hCE},
{8'hE5, 8'hE7, 8'hD0},
{8'hE0, 8'hE4, 8'hC9},
{8'hD0, 8'hD5, 8'hBA},
{8'hD3, 8'hD5, 8'hBB},
{8'hCA, 8'hB1, 8'h9A},
{8'hD9, 8'hBF, 8'hA9},
{8'hED, 8'hD7, 8'hC3},
{8'hFE, 8'hEF, 8'hE1},
{8'hFF, 8'hF7, 8'hF3},
{8'hFF, 8'hFA, 8'hFF},
{8'hD9, 8'hD2, 8'hE1},
{8'h11, 8'h0E, 8'h2A},
{8'h16, 8'h3E, 8'h84},
{8'h16, 8'h42, 8'h8C},
{8'h10, 8'h31, 8'h78},
{8'h0A, 8'h23, 8'h68},
{8'h12, 8'h29, 8'h6A},
{8'h13, 8'h24, 8'h5D},
{8'h05, 8'h0D, 8'h40},
{8'h00, 8'h00, 8'h2C},
{8'h02, 8'h03, 8'h24},
{8'h07, 8'h11, 8'h4E},
{8'h13, 8'h33, 8'h70},
{8'h06, 8'h24, 8'h44},
{8'h0A, 8'h32, 8'h56},
{8'h1E, 8'h38, 8'h7B},
{8'h42, 8'h4C, 8'h88},
{8'h6B, 8'h6A, 8'h7F},
{8'hA4, 8'h90, 8'h6E},
{8'hDB, 8'hD2, 8'h56},
{8'hE7, 8'hDA, 8'h4D},
{8'hF1, 8'hCD, 8'h97},
{8'hF4, 8'hC2, 8'hBC},
{8'hF5, 8'hC7, 8'h97},
{8'hF1, 8'hC7, 8'h79},
{8'hE5, 8'hCB, 8'h8E},
{8'hE1, 8'hD7, 8'h6C},
{8'hE9, 8'hD1, 8'h65},
{8'hC3, 8'hB4, 8'h72},
{8'h74, 8'h87, 8'h84},
{8'h24, 8'h44, 8'h68},
{8'h00, 8'h00, 8'h24},
{8'h02, 8'h00, 8'h17},
{8'h04, 8'h06, 8'h1E},
{8'h05, 8'h05, 8'h1A},
{8'h04, 8'h06, 8'h2C},
{8'h10, 8'h28, 8'h64},
{8'h1E, 8'h4B, 8'h9B},
{8'h1B, 8'h54, 8'hAE},
{8'h0B, 8'h44, 8'h9F},
{8'h0F, 8'h46, 8'h9F},
{8'h1B, 8'h55, 8'hAF},
{8'h19, 8'h52, 8'hC2},
{8'h20, 8'h50, 8'hBC},
{8'h37, 8'h55, 8'h8E},
{8'h84, 8'h8C, 8'h7D},
{8'hC1, 8'hB3, 8'h88},
{8'hFF, 8'hF3, 8'hDB},
{8'hFB, 8'hFB, 8'hE4},
{8'hF6, 8'hFD, 8'hD3},
{8'hFC, 8'hD7, 8'hB9},
{8'hF6, 8'hC2, 8'hA5},
{8'hFB, 8'hC2, 8'hA6},
{8'hFD, 8'hC2, 8'hA6},
{8'hFC, 8'hBC, 8'h9E},
{8'hF9, 8'hAF, 8'h8F},
{8'hF8, 8'hA6, 8'h89},
{8'hEE, 8'h96, 8'h77},
{8'hCA, 8'h97, 8'h70},
{8'hF1, 8'hD7, 8'hB2},
{8'hFC, 8'hF4, 8'hD1},
{8'hF2, 8'hF7, 8'hCC},
{8'hEF, 8'hF4, 8'hBE},
{8'hE9, 8'hED, 8'hB4},
{8'hF3, 8'hFC, 8'hC7},
{8'hD4, 8'hE3, 8'hB8},
{8'hAD, 8'hAD, 8'hA6},
{8'h88, 8'h87, 8'h84},
{8'h7E, 8'h7D, 8'h7B},
{8'h80, 8'h7F, 8'h7E},
{8'h7F, 8'h7D, 8'h7F},
{8'hFF, 8'hD7, 8'h00},
{8'h7F, 8'h7D, 8'h81},
{8'h7F, 8'h7D, 8'h82},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'h7F, 8'h7D, 8'h82},
{8'h7B, 8'h7A, 8'h87},
{8'h7C, 8'h80, 8'h6E},
{8'hCE, 8'hD8, 8'hA4},
{8'hE8, 8'hF6, 8'hB7},
{8'hE6, 8'hF4, 8'hBF},
{8'hE3, 8'hF2, 8'hC4},
{8'hE2, 8'hF4, 8'hBB},
{8'hE2, 8'hF5, 8'hAE},
{8'hE2, 8'hF2, 8'hA8},
{8'hE6, 8'hF5, 8'hB0},
{8'hE6, 8'hF2, 8'hB4},
{8'hE8, 8'hF1, 8'hBE},
{8'hE8, 8'hED, 8'hC4},
{8'hE3, 8'hE7, 8'hC4},
{8'hA1, 8'hA3, 8'h84},
{8'hA2, 8'hA2, 8'h88},
{8'hFC, 8'hF7, 8'hF9},
{8'hFA, 8'hF5, 8'hF6},
{8'hF6, 8'hF3, 8'hEC},
{8'hFB, 8'hFB, 8'hEC},
{8'hEB, 8'hEE, 8'hD8},
{8'hE7, 8'hEB, 8'hD2},
{8'hE7, 8'hEA, 8'hD2},
{8'hEA, 8'hEE, 8'hD6},
{8'hEC, 8'hE8, 8'hC4},
{8'hE0, 8'hDF, 8'hBC},
{8'hE6, 8'hEA, 8'hCF},
{8'hE8, 8'hF0, 8'hE3},
{8'hBB, 8'hCD, 8'hCB},
{8'h92, 8'hAB, 8'hB5},
{8'h42, 8'h61, 8'h77},
{8'h18, 8'h38, 8'h58},
{8'h1D, 8'h49, 8'h90},
{8'h1D, 8'h4C, 8'h98},
{8'h20, 8'h50, 8'h9E},
{8'h22, 8'h55, 8'hA4},
{8'h25, 8'h57, 8'hA5},
{8'h28, 8'h58, 8'hA3},
{8'h23, 8'h4F, 8'h98},
{8'h0F, 8'h30, 8'h73},
{8'h09, 8'h05, 8'h18},
{8'h06, 8'h01, 8'h2F},
{8'h07, 8'h0A, 8'h44},
{8'h04, 8'h10, 8'h37},
{8'h1D, 8'h29, 8'h47},
{8'h77, 8'h7C, 8'h8B},
{8'hB5, 8'hB8, 8'h89},
{8'hDA, 8'hDD, 8'h6C},
{8'hED, 8'hE0, 8'h9B},
{8'hF5, 8'hED, 8'hC4},
{8'hFE, 8'hFD, 8'hE1},
{8'hFB, 8'hFF, 8'hE7},
{8'hFA, 8'hFF, 8'hE7},
{8'hFC, 8'hFE, 8'hEA},
{8'hFD, 8'hFF, 8'hE6},
{8'hFC, 8'hFD, 8'hDE},
{8'hF1, 8'hE7, 8'hC6},
{8'hEC, 8'hCE, 8'h88},
{8'hEB, 8'hC7, 8'h63},
{8'hF4, 8'hDA, 8'h78},
{8'hCE, 8'hB6, 8'h64},
{8'h62, 8'h38, 8'h0C},
{8'h21, 8'h04, 8'h09},
{8'h07, 8'h00, 8'h31},
{8'h05, 8'h03, 8'h1F},
{8'h01, 8'h03, 8'h23},
{8'h03, 8'h10, 8'h41},
{8'h26, 8'h4C, 8'h92},
{8'h1C, 8'h4F, 8'hA9},
{8'h0F, 8'h48, 8'hA9},
{8'h1A, 8'h54, 8'hAF},
{8'h1B, 8'h57, 8'hAA},
{8'h19, 8'h5C, 8'h92},
{8'h57, 8'h70, 8'h7C},
{8'hCE, 8'hBC, 8'h8B},
{8'hFB, 8'hDA, 8'h89},
{8'hF9, 8'hE5, 8'hA8},
{8'hFE, 8'hFB, 8'hE4},
{8'hFD, 8'hF5, 8'hE1},
{8'hEF, 8'hDC, 8'hB5},
{8'hEC, 8'hBD, 8'h94},
{8'hEC, 8'hB3, 8'h8B},
{8'hEB, 8'hA5, 8'h7E},
{8'hF2, 8'hA0, 8'h7B},
{8'hF3, 8'hA0, 8'h79},
{8'hEB, 8'hA4, 8'h76},
{8'hD2, 8'hA3, 8'h6D},
{8'hD5, 8'hBC, 8'h80},
{8'hEE, 8'hE6, 8'hB0},
{8'hF2, 8'hF8, 8'hC6},
{8'hE8, 8'hFA, 8'hC9},
{8'hE5, 8'hF9, 8'hC3},
{8'hEC, 8'hF9, 8'hB8},
{8'hEF, 8'hF4, 8'hB4},
{8'hF1, 8'hF6, 8'hBE},
{8'hE7, 8'hF0, 8'hC4},
{8'hB5, 8'hB5, 8'hAE},
{8'h7C, 8'h7B, 8'h78},
{8'h83, 8'h82, 8'h80},
{8'h7B, 8'h7A, 8'h79},
{8'h7F, 8'h7D, 8'h7F},
{8'hFF, 8'hD7, 8'h00},
{8'h7F, 8'h7D, 8'h81},
{8'h7F, 8'h7D, 8'h82},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'h7E, 8'h7D, 8'h80},
{8'h7D, 8'h7D, 8'h83},
{8'h7A, 8'h7D, 8'h74},
{8'h94, 8'h9B, 8'h7F},
{8'hE7, 8'hF1, 8'hC8},
{8'hE4, 8'hF2, 8'hC0},
{8'hE3, 8'hF3, 8'hBC},
{8'hE2, 8'hF4, 8'hB7},
{8'hE3, 8'hF5, 8'hB4},
{8'hEA, 8'hFA, 8'hB4},
{8'hE5, 8'hF2, 8'hB3},
{8'hDF, 8'hE9, 8'hB4},
{8'hD8, 8'hE0, 8'hB5},
{8'hD9, 8'hDD, 8'hBC},
{8'hDC, 8'hDF, 8'hC3},
{8'hC6, 8'hC8, 8'hAE},
{8'hAE, 8'hAD, 8'h96},
{8'hF0, 8'hEC, 8'hE9},
{8'hF8, 8'hF5, 8'hF0},
{8'hF3, 8'hF1, 8'hE6},
{8'hF6, 8'hF6, 8'hE8},
{8'hF9, 8'hFB, 8'hEA},
{8'hFD, 8'hFE, 8'hEF},
{8'hFF, 8'hFF, 8'hFB},
{8'hFF, 8'hFF, 8'hFE},
{8'hE3, 8'hF0, 8'hF6},
{8'hA9, 8'hB9, 8'hC8},
{8'h60, 8'h79, 8'h97},
{8'h35, 8'h55, 8'h80},
{8'h14, 8'h44, 8'h7D},
{8'h0B, 8'h46, 8'h8D},
{8'h10, 8'h52, 8'hA3},
{8'h17, 8'h5D, 8'hB4},
{8'h15, 8'h56, 8'hB0},
{8'h14, 8'h57, 8'hB2},
{8'h10, 8'h56, 8'hB4},
{8'h0F, 8'h57, 8'hB5},
{8'h11, 8'h57, 8'hB6},
{8'h10, 8'h54, 8'hB0},
{8'h1B, 8'h5C, 8'hB5},
{8'h22, 8'h5D, 8'hAE},
{8'h14, 8'h23, 8'h32},
{8'h07, 8'h06, 8'h22},
{8'h09, 8'h00, 8'h22},
{8'h3D, 8'h25, 8'h27},
{8'hC1, 8'hA9, 8'h7A},
{8'hE6, 8'hDB, 8'h9B},
{8'hED, 8'hEC, 8'hB7},
{8'hF4, 8'hF6, 8'hD4},
{8'hFF, 8'hF6, 8'hEE},
{8'hFF, 8'hF8, 8'hF3},
{8'hFD, 8'hFB, 8'hF7},
{8'hF4, 8'hFF, 8'hF7},
{8'hED, 8'hFF, 8'hE3},
{8'hEF, 8'hFF, 8'hD1},
{8'hF6, 8'hFF, 8'hDB},
{8'hFB, 8'hFB, 8'hF2},
{8'hF5, 8'hFF, 8'hEA},
{8'hFB, 8'hFC, 8'hDB},
{8'hF9, 8'hEF, 8'hCB},
{8'hED, 8'hC7, 8'hA0},
{8'hF3, 8'h9F, 8'h63},
{8'hE8, 8'h76, 8'h32},
{8'h7F, 8'h35, 8'h19},
{8'h0C, 8'h00, 8'h10},
{8'h08, 8'h01, 8'h1C},
{8'h02, 8'h00, 8'h1A},
{8'h02, 8'h06, 8'h2B},
{8'h23, 8'h44, 8'h80},
{8'h16, 8'h42, 8'h9B},
{8'h14, 8'h48, 8'hAC},
{8'h1A, 8'h53, 8'hAE},
{8'h1F, 8'h59, 8'hA0},
{8'h69, 8'h85, 8'h66},
{8'hE0, 8'hDC, 8'h79},
{8'hFF, 8'hE8, 8'h6F},
{8'hF7, 8'hDC, 8'h94},
{8'hFC, 8'hF9, 8'hE6},
{8'hFC, 8'hFE, 8'hF5},
{8'hFA, 8'hE4, 8'hD3},
{8'hF9, 8'hD1, 8'hC1},
{8'hFC, 8'hEA, 8'hC2},
{8'hE6, 8'hCA, 8'h9E},
{8'hEE, 8'hC6, 8'h99},
{8'hF2, 8'hB8, 8'h8C},
{8'hE0, 8'h9E, 8'h72},
{8'hD3, 8'hAA, 8'h77},
{8'hEF, 8'hEC, 8'hAD},
{8'hE3, 8'hFB, 8'hB7},
{8'hE8, 8'hF5, 8'hBC},
{8'hE7, 8'hFC, 8'hC7},
{8'hDF, 8'hFD, 8'hC9},
{8'hE0, 8'hFB, 8'hC1},
{8'hEF, 8'hFB, 8'hBE},
{8'hEE, 8'hF2, 8'hB6},
{8'hF3, 8'hF8, 8'hC6},
{8'hE0, 8'hE8, 8'hC3},
{8'h8C, 8'h8C, 8'h86},
{8'h7C, 8'h7B, 8'h78},
{8'h83, 8'h82, 8'h80},
{8'h82, 8'h80, 8'h80},
{8'h80, 8'h7D, 8'h80},
{8'hFF, 8'hD7, 8'h00},
{8'h7F, 8'h7D, 8'h81},
{8'h7F, 8'h7D, 8'h82},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'h7F, 8'h7D, 8'h81},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'h7E, 8'h7D, 8'h7F},
{8'h7E, 8'h80, 8'h77},
{8'h85, 8'h86, 8'h87},
{8'h76, 8'h79, 8'h7C},
{8'hC3, 8'hCB, 8'hBC},
{8'hE6, 8'hF4, 8'hC8},
{8'hE3, 8'hF5, 8'hB5},
{8'hE2, 8'hF5, 8'hB4},
{8'hE3, 8'hF4, 8'hBC},
{8'hDF, 8'hEC, 8'hBA},
{8'hCD, 8'hD7, 8'hAD},
{8'hD7, 8'hDC, 8'hBE},
{8'hF2, 8'hF5, 8'hE2},
{8'hF8, 8'hF8, 8'hEB},
{8'hFE, 8'hFD, 8'hF2},
{8'hFB, 8'hF9, 8'hEF},
{8'hD3, 8'hCF, 8'hC4},
{8'hCA, 8'hC5, 8'hB8},
{8'hFF, 8'hFC, 8'hEE},
{8'hFD, 8'hF9, 8'hE8},
{8'hF7, 8'hF5, 8'hE4},
{8'hF7, 8'hF5, 8'hE7},
{8'hD1, 8'hD0, 8'hC8},
{8'hAA, 8'hA8, 8'hA6},
{8'h60, 8'h5E, 8'h63},
{8'h29, 8'h2A, 8'h48},
{8'h09, 8'h0D, 8'h36},
{8'h16, 8'h23, 8'h59},
{8'h1A, 8'h34, 8'h7A},
{8'h21, 8'h4B, 8'hA0},
{8'h1D, 8'h55, 8'hB7},
{8'h18, 8'h5A, 8'hC5},
{8'h14, 8'h5C, 8'hC9},
{8'h13, 8'h59, 8'hB8},
{8'h14, 8'h58, 8'hB5},
{8'h16, 8'h58, 8'hB3},
{8'h18, 8'h54, 8'hAB},
{8'h09, 8'h30, 8'h80},
{8'h03, 8'h21, 8'h6A},
{8'h0F, 8'h2F, 8'h71},
{8'h22, 8'h3F, 8'h82},
{8'h19, 8'h29, 8'h79},
{8'h00, 8'h01, 8'h0C},
{8'h0D, 8'h12, 8'h01},
{8'h9E, 8'h91, 8'h67},
{8'hFC, 8'hEA, 8'hCE},
{8'hFC, 8'hF5, 8'hE1},
{8'hFE, 8'hFC, 8'hE9},
{8'hF8, 8'hFA, 8'hEA},
{8'hFA, 8'hFD, 8'hCD},
{8'hFF, 8'hFE, 8'hD7},
{8'hFF, 8'hFC, 8'hDE},
{8'hF8, 8'hF7, 8'hD5},
{8'hFA, 8'hFE, 8'hD7},
{8'hFC, 8'hFF, 8'hDE},
{8'hFF, 8'hFA, 8'hE9},
{8'hFF, 8'hF6, 8'hF3},
{8'hF7, 8'hFD, 8'hF4},
{8'hF7, 8'hFB, 8'hE1},
{8'hFD, 8'hFF, 8'hE2},
{8'hF9, 8'hFE, 8'hE1},
{8'hFB, 8'hE9, 8'hB9},
{8'hF5, 8'hAC, 8'h6E},
{8'hD0, 8'h81, 8'h5B},
{8'h55, 8'h25, 8'h25},
{8'h0B, 8'h00, 8'h17},
{8'h03, 8'h00, 8'h14},
{8'h00, 8'h04, 8'h1E},
{8'h16, 8'h30, 8'h65},
{8'h13, 8'h35, 8'h8E},
{8'h1B, 8'h48, 8'hAE},
{8'h1A, 8'h4F, 8'hAA},
{8'h32, 8'h66, 8'hA3},
{8'hE5, 8'hD7, 8'h90},
{8'hF6, 8'hDE, 8'h7B},
{8'hF6, 8'hE3, 8'h8A},
{8'hFD, 8'hF7, 8'hC7},
{8'hF7, 8'hFB, 8'hF0},
{8'hF7, 8'hF9, 8'hF3},
{8'hFD, 8'hF3, 8'hE0},
{8'hFE, 8'hF2, 8'hD4},
{8'hF5, 8'hDC, 8'hC9},
{8'hF0, 8'hDE, 8'hC3},
{8'hFD, 8'hF4, 8'hD0},
{8'hFB, 8'hDD, 8'hB8},
{8'hF1, 8'hC0, 8'h9E},
{8'hD3, 8'hA3, 8'h81},
{8'hE1, 8'hD2, 8'hAA},
{8'hEE, 8'hF8, 8'hCB},
{8'hF6, 8'hF5, 8'hC5},
{8'hE9, 8'hF2, 8'hC5},
{8'hE4, 8'hF7, 8'hCA},
{8'hE9, 8'hFB, 8'hC9},
{8'hE8, 8'hF2, 8'hB9},
{8'hF3, 8'hF7, 8'hC2},
{8'hF1, 8'hFA, 8'hD2},
{8'h9D, 8'hAA, 8'h90},
{8'h7B, 8'h7C, 8'h76},
{8'h7C, 8'h7B, 8'h78},
{8'h84, 8'h83, 8'h80},
{8'h7B, 8'h7A, 8'h79},
{8'h7E, 8'h7C, 8'h7E},
{8'hFF, 8'hD7, 8'h00},
{8'h7F, 8'h7D, 8'h81},
{8'h7F, 8'h7D, 8'h82},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'h81, 8'h7C, 8'h7F},
{8'h81, 8'h7C, 8'h7F},
{8'h80, 8'h7C, 8'h7F},
{8'h80, 8'h7C, 8'h7F},
{8'h80, 8'h7D, 8'h7F},
{8'h7F, 8'h7D, 8'h7F},
{8'h7F, 8'h7D, 8'h7F},
{8'h7F, 8'h7D, 8'h7F},
{8'h7D, 8'h7E, 8'h80},
{8'h7E, 8'h7E, 8'h7F},
{8'h7E, 8'h7E, 8'h7F},
{8'h7F, 8'h7E, 8'h7E},
{8'h7F, 8'h7E, 8'h7E},
{8'h7F, 8'h7E, 8'h7E},
{8'h7E, 8'h7E, 8'h7E},
{8'h7E, 8'h7E, 8'h7E},
{8'h82, 8'h7D, 8'h7A},
{8'h81, 8'h7C, 8'h7E},
{8'h80, 8'h7C, 8'h82},
{8'h7F, 8'h7D, 8'h84},
{8'h80, 8'h7E, 8'h82},
{8'h80, 8'h7D, 8'h7F},
{8'h81, 8'h7C, 8'h7D},
{8'h82, 8'h7C, 8'h7E},
{8'h7B, 8'h7C, 8'h7B},
{8'h7E, 8'h7C, 8'h87},
{8'h7D, 8'h7A, 8'h89},
{8'h92, 8'h93, 8'h8F},
{8'hE6, 8'hEC, 8'hC5},
{8'hE7, 8'hF3, 8'hB3},
{8'hE6, 8'hF6, 8'hB4},
{8'hDE, 8'hED, 8'hB4},
{8'hD3, 8'hDA, 8'hAB},
{8'hE7, 8'hEC, 8'hC7},
{8'hFB, 8'hFE, 8'hE8},
{8'hFF, 8'hFF, 8'hFD},
{8'hF4, 8'hFA, 8'hFC},
{8'hE9, 8'hF2, 8'hF9},
{8'hDD, 8'hE8, 8'hEF},
{8'hD3, 8'hE0, 8'hE6},
{8'hB7, 8'hBD, 8'hC9},
{8'hB0, 8'hB6, 8'hC3},
{8'h9A, 8'hA3, 8'hB1},
{8'h66, 8'h73, 8'h84},
{8'h34, 8'h45, 8'h5D},
{8'h12, 8'h24, 8'h40},
{8'h00, 8'h0F, 8'h2F},
{8'h00, 8'h0B, 8'h2F},
{8'h0E, 8'h0C, 8'h27},
{8'h09, 8'h0A, 8'h24},
{8'h02, 8'h05, 8'h23},
{8'h00, 8'h04, 8'h28},
{8'h03, 8'h0C, 8'h39},
{8'h07, 8'h1D, 8'h53},
{8'h12, 8'h35, 8'h74},
{8'h1F, 8'h47, 8'h8C},
{8'h22, 8'h54, 8'hA7},
{8'h21, 8'h55, 8'hA6},
{8'h23, 8'h56, 8'hA4},
{8'h25, 8'h52, 8'hA0},
{8'h22, 8'h43, 8'h8F},
{8'h0A, 8'h18, 8'h59},
{8'h00, 8'h00, 8'h2D},
{8'h04, 8'h01, 8'h26},
{8'h07, 8'h11, 8'h3A},
{8'h34, 8'h3A, 8'h51},
{8'h9F, 8'hA7, 8'hB4},
{8'hE8, 8'hEC, 8'hF6},
{8'hF2, 8'hF5, 8'hE5},
{8'hFA, 8'hFD, 8'hCA},
{8'hFE, 8'hFE, 8'hD3},
{8'hFD, 8'hFA, 8'hEC},
{8'hF1, 8'hFF, 8'hCE},
{8'hF9, 8'hFD, 8'hE2},
{8'hEE, 8'hE7, 8'hDE},
{8'hF2, 8'hEA, 8'hDA},
{8'hF8, 8'hF5, 8'hD5},
{8'hF9, 8'hF6, 8'hD8},
{8'hF8, 8'hF4, 8'hDD},
{8'hF8, 8'hF2, 8'hE1},
{8'hF8, 8'hF1, 8'hE9},
{8'hFE, 8'hF8, 8'hDC},
{8'hFC, 8'hFE, 8'hDB},
{8'hE7, 8'hFE, 8'hE8},
{8'hEA, 8'hFF, 8'hEF},
{8'hFB, 8'hF2, 8'hC7},
{8'hF9, 8'hC5, 8'h8B},
{8'hDD, 8'h9B, 8'h65},
{8'h3A, 8'h22, 8'h2D},
{8'h06, 8'h01, 8'h13},
{8'h01, 8'h03, 8'h1E},
{8'h03, 8'h0A, 8'h33},
{8'h0E, 8'h1F, 8'h61},
{8'h26, 8'h47, 8'hA0},
{8'h1D, 8'h4F, 8'hAB},
{8'h2F, 8'h64, 8'hA6},
{8'hEF, 8'hCE, 8'h8A},
{8'hF7, 8'hDA, 8'hA6},
{8'hF9, 8'hF8, 8'hD8},
{8'hF6, 8'hFE, 8'hDE},
{8'hF8, 8'hF8, 8'hE0},
{8'hFE, 8'hF3, 8'hE6},
{8'hFB, 8'hE3, 8'hC5},
{8'hEA, 8'hCF, 8'h95},
{8'hF2, 8'hD0, 8'hC2},
{8'hFF, 8'hF2, 8'hE4},
{8'hFF, 8'hF8, 8'hE2},
{8'hFD, 8'hF9, 8'hE2},
{8'hF9, 8'hE8, 8'hD3},
{8'hF9, 8'hD1, 8'hBF},
{8'hE3, 8'hC1, 8'hAC},
{8'hFA, 8'hE4, 8'hCB},
{8'hF8, 8'hEE, 8'hC2},
{8'hEE, 8'hEE, 8'hC3},
{8'hC7, 8'hCE, 8'hA6},
{8'hB8, 8'hC1, 8'h96},
{8'hE0, 8'hE6, 8'hB8},
{8'hE2, 8'hE7, 8'hBF},
{8'hB7, 8'hC0, 8'hA2},
{8'hB5, 8'hC3, 8'hB0},
{8'h7C, 8'h7C, 8'h79},
{8'h84, 8'h82, 8'h81},
{8'h7C, 8'h7A, 8'h7A},
{8'h7C, 8'h7B, 8'h7C},
{8'h7E, 8'h7C, 8'h7F},
{8'h7F, 8'h7D, 8'h7F},
{8'h7F, 8'h7D, 8'h7F},
{8'h7F, 8'h7E, 8'h7F},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'h84, 8'h7B, 8'h7F},
{8'h84, 8'h7B, 8'h7F},
{8'h83, 8'h7C, 8'h7F},
{8'h82, 8'h7C, 8'h7F},
{8'h81, 8'h7C, 8'h7F},
{8'h7F, 8'h7D, 8'h7F},
{8'h7F, 8'h7D, 8'h7F},
{8'h7E, 8'h7E, 8'h7F},
{8'h7B, 8'h7F, 8'h80},
{8'h7C, 8'h7F, 8'h7E},
{8'h7E, 8'h7F, 8'h7B},
{8'h7F, 8'h7E, 8'h7A},
{8'h7F, 8'h7E, 8'h7A},
{8'h7E, 8'h7F, 8'h7A},
{8'h7D, 8'h7F, 8'h7C},
{8'h7D, 8'h7F, 8'h7C},
{8'h84, 8'h7D, 8'h76},
{8'h82, 8'h7C, 8'h7D},
{8'h7E, 8'h7D, 8'h84},
{8'h7A, 8'h7F, 8'h81},
{8'h7A, 8'h7F, 8'h79},
{8'h80, 8'h80, 8'h7D},
{8'h85, 8'h7C, 8'h88},
{8'h83, 8'h75, 8'h8F},
{8'h77, 8'h75, 8'h93},
{8'h7F, 8'h7C, 8'h90},
{8'h82, 8'h7E, 8'h7D},
{8'h7F, 8'h7C, 8'h66},
{8'hCB, 8'hCD, 8'hA3},
{8'hF1, 8'hFA, 8'hC1},
{8'hE5, 8'hF7, 8'hB4},
{8'hC4, 8'hDD, 8'h97},
{8'hBE, 8'hCF, 8'hC1},
{8'h9E, 8'hB0, 8'hB2},
{8'h86, 8'h9C, 8'hB2},
{8'h52, 8'h6B, 8'h97},
{8'h3C, 8'h58, 8'h92},
{8'h30, 8'h58, 8'h99},
{8'h24, 8'h55, 8'h96},
{8'h1F, 8'h54, 8'h95},
{8'h21, 8'h48, 8'hA4},
{8'h12, 8'h3D, 8'h9E},
{8'h0D, 8'h3F, 8'hA2},
{8'h11, 8'h4D, 8'hB2},
{8'h0F, 8'h51, 8'hB6},
{8'h0F, 8'h55, 8'hB9},
{8'h0F, 8'h55, 8'hB7},
{8'h0F, 8'h53, 8'hB0},
{8'h14, 8'h52, 8'hA2},
{8'h13, 8'h4D, 8'h9E},
{8'h12, 8'h46, 8'h98},
{8'h16, 8'h41, 8'h90},
{8'h16, 8'h3A, 8'h82},
{8'h0E, 8'h2E, 8'h6B},
{8'h08, 8'h23, 8'h55},
{8'h0D, 8'h23, 8'h50},
{8'h10, 8'h27, 8'h74},
{8'h18, 8'h3C, 8'h85},
{8'h17, 8'h50, 8'h98},
{8'h18, 8'h57, 8'hB1},
{8'h1C, 8'h54, 8'hC0},
{8'h28, 8'h50, 8'hB4},
{8'h19, 8'h30, 8'h6E},
{8'h15, 8'h22, 8'h3C},
{8'h92, 8'h91, 8'h96},
{8'hF4, 8'hF3, 8'hF5},
{8'hFF, 8'hFF, 8'hFF},
{8'hF6, 8'hFB, 8'hF6},
{8'hED, 8'hF2, 8'hE5},
{8'hED, 8'hEE, 8'hDE},
{8'hFA, 8'hF9, 8'hE6},
{8'hFF, 8'hFC, 8'hE5},
{8'hFF, 8'hFA, 8'hDF},
{8'hEE, 8'hE5, 8'hCC},
{8'hF2, 8'hEB, 8'hD5},
{8'hF4, 8'hF0, 8'hE0},
{8'hF9, 8'hF5, 8'hEB},
{8'hF9, 8'hF6, 8'hF1},
{8'hF8, 8'hF6, 8'hF5},
{8'hF8, 8'hF6, 8'hF8},
{8'hF7, 8'hF6, 8'hF8},
{8'hF8, 8'hF1, 8'hE8},
{8'hF9, 8'hF0, 8'hD8},
{8'hF9, 8'hF6, 8'hDD},
{8'hF4, 8'hFA, 8'hE9},
{8'hFD, 8'hFF, 8'hEB},
{8'hFA, 8'hE2, 8'hBC},
{8'hFF, 8'hC2, 8'h8B},
{8'h6E, 8'h54, 8'h3D},
{8'h04, 8'h00, 8'h11},
{8'h01, 8'h01, 8'h2C},
{8'h00, 8'h01, 8'h11},
{8'h04, 8'h04, 8'h0D},
{8'h30, 8'h3B, 8'h70},
{8'h24, 8'h4E, 8'hAD},
{8'h18, 8'h55, 8'hAD},
{8'hC5, 8'h9C, 8'h6A},
{8'hFD, 8'hED, 8'hBE},
{8'hF2, 8'hFF, 8'hE8},
{8'hEF, 8'hFF, 8'hF2},
{8'hFD, 8'hF7, 8'hE5},
{8'hFE, 8'hD8, 8'hB8},
{8'hF5, 8'hB2, 8'h84},
{8'hFA, 8'hBD, 8'h87},
{8'hFB, 8'hF0, 8'hCE},
{8'hFF, 8'hFA, 8'hE1},
{8'hFB, 8'hF7, 8'hE5},
{8'hF6, 8'hFD, 8'hEE},
{8'hF0, 8'hFF, 8'hED},
{8'hF3, 8'hFC, 8'hE4},
{8'hE4, 8'hD9, 8'hBC},
{8'hE9, 8'hD0, 8'hAE},
{8'hF0, 8'hFC, 8'hC2},
{8'hEC, 8'hF8, 8'hC1},
{8'hEB, 8'hF4, 8'hC6},
{8'hED, 8'hF5, 8'hD0},
{8'hD8, 8'hDD, 8'hC0},
{8'h85, 8'h89, 8'h73},
{8'h78, 8'h7A, 8'h67},
{8'hCE, 8'hCE, 8'hBE},
{8'h93, 8'h92, 8'h90},
{8'h81, 8'h7E, 8'h81},
{8'h7E, 8'h7C, 8'h81},
{8'h7E, 8'h7B, 8'h82},
{8'h7E, 8'h7C, 8'h81},
{8'h7F, 8'h7D, 8'h7E},
{8'h7F, 8'h7E, 8'h79},
{8'h7F, 8'h7F, 8'h77},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'h7E, 8'h7E, 8'h80},
{8'h7E, 8'h7E, 8'h80},
{8'h7E, 8'h7E, 8'h80},
{8'h7E, 8'h7E, 8'h80},
{8'h82, 8'h7C, 8'h7F},
{8'h82, 8'h7C, 8'h7F},
{8'h83, 8'h7C, 8'h7E},
{8'h83, 8'h7C, 8'h7E},
{8'h82, 8'h7C, 8'h7F},
{8'h82, 8'h7C, 8'h80},
{8'h81, 8'h7C, 8'h81},
{8'h7F, 8'h7D, 8'h83},
{8'h78, 8'h80, 8'h87},
{8'h77, 8'h7F, 8'h8A},
{8'h77, 8'h80, 8'h88},
{8'h77, 8'h81, 8'h7F},
{8'h7A, 8'h85, 8'h77},
{8'h79, 8'h84, 8'h78},
{8'h78, 8'h7F, 8'h85},
{8'h77, 8'h7B, 8'h8F},
{8'h7B, 8'h80, 8'h79},
{8'h7F, 8'h83, 8'h79},
{8'h7D, 8'h81, 8'h79},
{8'h7B, 8'h82, 8'h7E},
{8'h88, 8'h96, 8'h97},
{8'hB2, 8'hC8, 8'hD1},
{8'h70, 8'h8E, 8'hA0},
{8'h38, 8'h5E, 8'h77},
{8'h1B, 8'h59, 8'h9B},
{8'h0F, 8'h4E, 8'h9B},
{8'h12, 8'h4E, 8'hA7},
{8'h10, 8'h4A, 8'hAF},
{8'h14, 8'h4D, 8'hB7},
{8'h16, 8'h4F, 8'hB8},
{8'h19, 8'h52, 8'hB7},
{8'h1B, 8'h55, 8'hB4},
{8'h19, 8'h56, 8'hB1},
{8'h1A, 8'h5A, 8'hB5},
{8'h18, 8'h5A, 8'hB7},
{8'h13, 8'h58, 8'hB4},
{8'h16, 8'h5A, 8'hB3},
{8'h17, 8'h59, 8'hAD},
{8'h1A, 8'h57, 8'hA7},
{8'h1C, 8'h57, 8'hA7},
{8'h15, 8'h53, 8'hBA},
{8'h15, 8'h53, 8'hBC},
{8'h15, 8'h55, 8'hBC},
{8'h15, 8'h56, 8'hBD},
{8'h16, 8'h57, 8'hBE},
{8'h1B, 8'h5D, 8'hC5},
{8'h18, 8'h5B, 8'hC5},
{8'h10, 8'h51, 8'hBC},
{8'h18, 8'h4B, 8'hA4},
{8'h0E, 8'h43, 8'h94},
{8'h07, 8'h45, 8'h92},
{8'h08, 8'h4E, 8'hA3},
{8'h11, 8'h50, 8'hAC},
{8'h1D, 8'h4B, 8'h99},
{8'h43, 8'h61, 8'h8A},
{8'hC0, 8'hCF, 8'hD8},
{8'hFF, 8'hFF, 8'hFF},
{8'hFE, 8'hFF, 8'hFF},
{8'hF6, 8'hFA, 8'hF6},
{8'hFA, 8'hFE, 8'hF8},
{8'hFD, 8'hFF, 8'hF7},
{8'hF8, 8'hFA, 8'hED},
{8'hF1, 8'hEE, 8'hDF},
{8'hF4, 8'hF0, 8'hE0},
{8'hE4, 8'hE1, 8'hCE},
{8'hE8, 8'hE3, 8'hD1},
{8'hFC, 8'hFB, 8'hEB},
{8'hFD, 8'hFD, 8'hF1},
{8'hFF, 8'hFF, 8'hF7},
{8'hFF, 8'hFF, 8'hFA},
{8'hFF, 8'hFF, 8'hFD},
{8'hFF, 8'hFF, 8'hFE},
{8'hFD, 8'hFF, 8'hFF},
{8'hFE, 8'hFD, 8'hF6},
{8'hFE, 8'hFB, 8'hE8},
{8'hF6, 8'hF6, 8'hE3},
{8'hEF, 8'hF4, 8'hE5},
{8'hFB, 8'hF7, 8'hE8},
{8'hFF, 8'hF1, 8'hD5},
{8'hFD, 8'hCD, 8'hA4},
{8'h6B, 8'h54, 8'h44},
{8'h00, 8'h00, 8'h0F},
{8'h04, 8'h01, 8'h2C},
{8'h02, 8'h04, 8'h18},
{8'h06, 8'h08, 8'h15},
{8'h07, 8'h0B, 8'h39},
{8'h0B, 8'h27, 8'h79},
{8'h15, 8'h4D, 8'h9D},
{8'h86, 8'h78, 8'h6E},
{8'hFE, 8'hFA, 8'hE7},
{8'hF9, 8'hFD, 8'hE5},
{8'hFD, 8'hFC, 8'hE1},
{8'hFE, 8'hEF, 8'hCF},
{8'hEC, 8'hC2, 8'hA2},
{8'hEB, 8'hC3, 8'hA3},
{8'hFB, 8'hE6, 8'hC7},
{8'hFF, 8'hFC, 8'hE3},
{8'hFC, 8'hF6, 8'hDF},
{8'hFB, 8'hF3, 8'hDE},
{8'hFC, 8'hFA, 8'hE4},
{8'hFA, 8'hFA, 8'hE1},
{8'hF0, 8'hEF, 8'hD3},
{8'hF6, 8'hEE, 8'hD3},
{8'hE1, 8'hD0, 8'hB3},
{8'hE5, 8'hEC, 8'hBA},
{8'hED, 8'hF7, 8'hC5},
{8'hE9, 8'hF1, 8'hC4},
{8'hF0, 8'hF7, 8'hCF},
{8'hEA, 8'hEF, 8'hCC},
{8'hB7, 8'hBB, 8'h9D},
{8'h80, 8'h84, 8'h66},
{8'hD3, 8'hD5, 8'hBC},
{8'hAF, 8'hAE, 8'hA7},
{8'h78, 8'h77, 8'h74},
{8'h80, 8'h7E, 8'h80},
{8'h81, 8'h7F, 8'h84},
{8'h7F, 8'h7C, 8'h82},
{8'h7F, 8'h7D, 8'h81},
{8'h7F, 8'h7E, 8'h7D},
{8'h7F, 8'h7E, 8'h7C},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'h7A, 8'h80, 8'h80},
{8'h7B, 8'h80, 8'h80},
{8'h7B, 8'h7F, 8'h80},
{8'h7C, 8'h7E, 8'h80},
{8'h7D, 8'h7E, 8'h80},
{8'h7E, 8'h7E, 8'h80},
{8'h7E, 8'h7D, 8'h80},
{8'h80, 8'h7D, 8'h80},
{8'h86, 8'h7A, 8'h7E},
{8'h86, 8'h7A, 8'h7F},
{8'h85, 8'h7B, 8'h81},
{8'h83, 8'h7B, 8'h83},
{8'h82, 8'h7B, 8'h83},
{8'h81, 8'h7B, 8'h84},
{8'h81, 8'h7B, 8'h84},
{8'h80, 8'h7C, 8'h83},
{8'h7B, 8'h81, 8'h77},
{8'h7C, 8'h7E, 8'h84},
{8'h81, 8'h79, 8'h92},
{8'h83, 8'h78, 8'h91},
{8'h81, 8'h7B, 8'h80},
{8'h80, 8'h81, 8'h70},
{8'h7F, 8'h88, 8'h69},
{8'h7F, 8'h8A, 8'h69},
{8'h86, 8'h84, 8'h74},
{8'h81, 8'h7E, 8'h78},
{8'h74, 8'h72, 8'h7A},
{8'h53, 8'h53, 8'h6E},
{8'h2E, 8'h32, 8'h64},
{8'h1F, 8'h27, 8'h6F},
{8'h0F, 8'h1B, 8'h76},
{8'h0C, 8'h1D, 8'h7E},
{8'h04, 8'h2E, 8'h75},
{8'h0E, 8'h3B, 8'h86},
{8'h16, 8'h46, 8'h9E},
{8'h1B, 8'h50, 8'hB2},
{8'h1A, 8'h53, 8'hBB},
{8'h16, 8'h55, 8'hBC},
{8'h14, 8'h56, 8'hBD},
{8'h14, 8'h57, 8'hBA},
{8'h0F, 8'h5B, 8'hB4},
{8'h0A, 8'h57, 8'hB1},
{8'h0A, 8'h57, 8'hB1},
{8'h0F, 8'h5B, 8'hB5},
{8'h12, 8'h5A, 8'hB1},
{8'h0E, 8'h4F, 8'hA2},
{8'h14, 8'h4E, 8'h9D},
{8'h1F, 8'h57, 8'hA3},
{8'h1C, 8'h51, 8'hA9},
{8'h1C, 8'h53, 8'hAB},
{8'h1B, 8'h57, 8'hAF},
{8'h1A, 8'h58, 8'hB2},
{8'h17, 8'h59, 8'hB7},
{8'h14, 8'h58, 8'hBD},
{8'h11, 8'h58, 8'hC3},
{8'h10, 8'h57, 8'hC5},
{8'h18, 8'h57, 8'hB6},
{8'h16, 8'h5B, 8'hB3},
{8'h12, 8'h5D, 8'hAF},
{8'h0F, 8'h57, 8'hA6},
{8'h0F, 8'h4C, 8'h95},
{8'h43, 8'h6B, 8'h9A},
{8'hD2, 8'hE6, 8'hEB},
{8'hFA, 8'hFF, 8'hFD},
{8'hFC, 8'hFC, 8'hF7},
{8'hF9, 8'hFB, 8'hF5},
{8'hF9, 8'hFC, 8'hF6},
{8'hFB, 8'hFE, 8'hF9},
{8'hFC, 8'hFE, 8'hF8},
{8'hFD, 8'hFE, 8'hF7},
{8'hFA, 8'hF7, 8'hF0},
{8'hD2, 8'hCA, 8'hC4},
{8'hDF, 8'hDE, 8'hD7},
{8'hFD, 8'hFD, 8'hF8},
{8'hFC, 8'hFC, 8'hF6},
{8'hFA, 8'hFA, 8'hF5},
{8'hFD, 8'hFE, 8'hF9},
{8'hFD, 8'hFE, 8'hFA},
{8'hFD, 8'hFF, 8'hFA},
{8'hFB, 8'hFF, 8'hFB},
{8'hF9, 8'hFF, 8'hFF},
{8'hFD, 8'hFD, 8'hFA},
{8'hFE, 8'hFE, 8'hF4},
{8'hFD, 8'hFE, 8'hF3},
{8'hFD, 8'hFF, 8'hF7},
{8'hF9, 8'hF0, 8'hE7},
{8'hFC, 8'hE1, 8'hD3},
{8'hF0, 8'hC9, 8'hB2},
{8'h54, 8'h44, 8'h3C},
{8'h01, 8'h00, 8'h11},
{8'h07, 8'h02, 8'h2A},
{8'h02, 8'h02, 8'h1C},
{8'h06, 8'h06, 8'h19},
{8'h00, 8'h03, 8'h2A},
{8'h1A, 8'h36, 8'h76},
{8'h2C, 8'h56, 8'h9A},
{8'h68, 8'h70, 8'h8A},
{8'hEF, 8'hF1, 8'hF6},
{8'hFF, 8'hFA, 8'hEA},
{8'hFF, 8'hF8, 8'hD8},
{8'hFC, 8'hE6, 8'hC4},
{8'hF0, 8'hD1, 8'hB7},
{8'hF4, 8'hE8, 8'hD6},
{8'hFA, 8'hFE, 8'hF1},
{8'hFA, 8'hF9, 8'hE9},
{8'hFB, 8'hF4, 8'hE0},
{8'hFF, 8'hF9, 8'hE0},
{8'hFF, 8'hF9, 8'hDD},
{8'hF8, 8'hE5, 8'hC8},
{8'hFD, 8'hEF, 8'hD4},
{8'hFF, 8'hFA, 8'hE2},
{8'hEE, 8'hEA, 8'hD4},
{8'hD9, 8'hDD, 8'hB6},
{8'hF0, 8'hF6, 8'hCB},
{8'hED, 8'hF3, 8'hC7},
{8'hEF, 8'hF6, 8'hCA},
{8'hED, 8'hF2, 8'hC8},
{8'hED, 8'hF3, 8'hCA},
{8'hD6, 8'hDD, 8'hB3},
{8'hF0, 8'hF6, 8'hD0},
{8'hD5, 8'hD7, 8'hC8},
{8'h81, 8'h80, 8'h78},
{8'h83, 8'h81, 8'h7F},
{8'h80, 8'h7E, 8'h82},
{8'h7F, 8'h7B, 8'h83},
{8'h7F, 8'h7C, 8'h83},
{8'h7F, 8'h7D, 8'h82},
{8'h7F, 8'h7D, 8'h82},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'h79, 8'h7F, 8'h7D},
{8'h79, 8'h7F, 8'h7D},
{8'h7C, 8'h80, 8'h7E},
{8'h7D, 8'h7E, 8'h7D},
{8'h7E, 8'h7E, 8'h7E},
{8'h80, 8'h7E, 8'h7E},
{8'h82, 8'h7F, 8'h80},
{8'h80, 8'h7C, 8'h7D},
{8'h82, 8'h7A, 8'h7B},
{8'h82, 8'h7C, 8'h7F},
{8'h7D, 8'h7B, 8'h81},
{8'h7D, 8'h7E, 8'h84},
{8'h7D, 8'h7E, 8'h86},
{8'h7D, 8'h7E, 8'h84},
{8'h7D, 8'h7C, 8'h80},
{8'h80, 8'h7B, 8'h7D},
{8'h82, 8'h81, 8'h6B},
{8'h85, 8'h7F, 8'h73},
{8'h84, 8'h79, 8'h7A},
{8'h87, 8'h7A, 8'h7D},
{8'h85, 8'h7C, 8'h7D},
{8'h85, 8'h81, 8'h88},
{8'h63, 8'h65, 8'h7B},
{8'h4C, 8'h50, 8'h76},
{8'h51, 8'h55, 8'h84},
{8'h3C, 8'h41, 8'h6C},
{8'h14, 8'h15, 8'h39},
{8'h00, 8'h00, 8'h1B},
{8'h00, 8'h02, 8'h17},
{8'h00, 8'h03, 8'h10},
{8'h00, 8'h05, 8'h0E},
{8'h00, 8'h06, 8'h0D},
{8'h04, 8'h00, 8'h13},
{8'h01, 8'h00, 8'h1C},
{8'h03, 8'h08, 8'h32},
{8'h07, 8'h18, 8'h50},
{8'h13, 8'h30, 8'h71},
{8'h12, 8'h3D, 8'h87},
{8'h15, 8'h4F, 8'h9B},
{8'h1A, 8'h5B, 8'hA8},
{8'h16, 8'h5B, 8'hAE},
{8'h15, 8'h5B, 8'hB1},
{8'h12, 8'h5A, 8'hB4},
{8'h0F, 8'h57, 8'hB5},
{8'h0E, 8'h57, 8'hB5},
{8'h11, 8'h56, 8'hB4},
{8'h07, 8'h45, 8'hA1},
{8'h08, 8'h35, 8'h8D},
{8'h0D, 8'h2C, 8'h66},
{8'h05, 8'h2A, 8'h67},
{8'h05, 8'h2C, 8'h70},
{8'h0B, 8'h30, 8'h7B},
{8'h0E, 8'h35, 8'h81},
{8'h17, 8'h43, 8'h8B},
{8'h20, 8'h4B, 8'h8E},
{8'h25, 8'h51, 8'h92},
{8'h1A, 8'h50, 8'hA8},
{8'h1B, 8'h54, 8'hAB},
{8'h1A, 8'h54, 8'hA5},
{8'h1C, 8'h52, 8'h98},
{8'h3D, 8'h66, 8'h9A},
{8'hD0, 8'hE5, 8'hEF},
{8'hFF, 8'hFF, 8'hFF},
{8'hFE, 8'hFA, 8'hF0},
{8'hFE, 8'hFC, 8'hF4},
{8'hFE, 8'hFE, 8'hF7},
{8'hFD, 8'hFD, 8'hF7},
{8'hFC, 8'hFE, 8'hF8},
{8'hFD, 8'hFD, 8'hF8},
{8'hFF, 8'hFF, 8'hFD},
{8'hE9, 8'hE0, 8'hE1},
{8'hD0, 8'hC4, 8'hC7},
{8'hFA, 8'hF9, 8'hFA},
{8'hFB, 8'hFB, 8'hFC},
{8'hFC, 8'hFB, 8'hFC},
{8'hFE, 8'hFE, 8'hFE},
{8'hFD, 8'hFE, 8'hFC},
{8'hFD, 8'hFE, 8'hFB},
{8'hFD, 8'hFE, 8'hFA},
{8'hFD, 8'hFF, 8'hFA},
{8'hFA, 8'hFE, 8'hFF},
{8'hFB, 8'hFE, 8'hFF},
{8'hFD, 8'hFE, 8'hFD},
{8'hFF, 8'hFF, 8'hFC},
{8'hFF, 8'hFA, 8'hF8},
{8'hFF, 8'hFC, 8'hFA},
{8'hF6, 8'hDF, 8'hDD},
{8'hC6, 8'hA3, 8'hA1},
{8'h2E, 8'h27, 8'h2C},
{8'h05, 8'h01, 8'h15},
{8'h06, 8'h01, 8'h23},
{8'h04, 8'h00, 8'h21},
{8'h03, 8'h06, 8'h1F},
{8'h01, 8'h03, 8'h1E},
{8'h04, 8'h11, 8'h39},
{8'h1A, 8'h2E, 8'h5F},
{8'h55, 8'h59, 8'h7F},
{8'hE1, 8'hDE, 8'hEE},
{8'hFF, 8'hF8, 8'hF0},
{8'hFE, 8'hF5, 8'hE0},
{8'hFD, 8'hF2, 8'hDE},
{8'hFF, 8'hFA, 8'hEA},
{8'hFA, 8'hF9, 8'hE9},
{8'hF4, 8'hF9, 8'hE7},
{8'hFE, 8'hFD, 8'hF0},
{8'hFF, 8'hFA, 8'hE8},
{8'hFF, 8'hF6, 8'hDA},
{8'hFB, 8'hDF, 8'hC0},
{8'hEA, 8'hBC, 8'h9F},
{8'hFE, 8'hE2, 8'hCA},
{8'hFE, 8'hF6, 8'hE0},
{8'hFA, 8'hFD, 8'hE9},
{8'hDB, 8'hDD, 8'hBE},
{8'hCE, 8'hCF, 8'hAC},
{8'hD9, 8'hDB, 8'hB2},
{8'hD7, 8'hDB, 8'hAC},
{8'hE5, 8'hEB, 8'hBA},
{8'hEF, 8'hF7, 8'hC4},
{8'hEF, 8'hF6, 8'hC5},
{8'hF1, 8'hF8, 8'hCB},
{8'hC4, 8'hC6, 8'hB4},
{8'h79, 8'h79, 8'h6E},
{8'h7C, 8'h7B, 8'h78},
{8'h83, 8'h81, 8'h84},
{8'h80, 8'h7D, 8'h85},
{8'h7F, 8'h7C, 8'h85},
{8'h7F, 8'h7C, 8'h85},
{8'h7F, 8'h7C, 8'h83},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'h80, 8'h7D, 8'h80},
{8'h7F, 8'h7A, 8'h78},
{8'h7C, 8'h78, 8'h74},
{8'h82, 8'h7C, 8'h79},
{8'h80, 8'h7A, 8'h77},
{8'h7F, 8'h7A, 8'h77},
{8'h7D, 8'h77, 8'h73},
{8'h7A, 8'h74, 8'h71},
{8'h81, 8'h79, 8'h77},
{8'h7A, 8'h79, 8'h73},
{8'h7C, 8'h7F, 8'h7B},
{8'h7C, 8'h83, 8'h82},
{8'h77, 8'h80, 8'h81},
{8'h75, 8'h7C, 8'h7C},
{8'h7E, 8'h80, 8'h7C},
{8'h82, 8'h7F, 8'h75},
{8'h82, 8'h7B, 8'h71},
{8'h79, 8'h7C, 8'h89},
{8'h76, 8'h7E, 8'h8A},
{8'h67, 8'h78, 8'h7C},
{8'h53, 8'h6D, 8'h6B},
{8'h4D, 8'h6B, 8'h73},
{8'h38, 8'h57, 8'h85},
{8'h27, 8'h40, 8'hA6},
{8'h26, 8'h3E, 8'hC6},
{8'h14, 8'h46, 8'h9C},
{8'h17, 8'h4A, 8'h99},
{8'h14, 8'h42, 8'h8E},
{8'h14, 8'h3B, 8'h82},
{8'h0C, 8'h2E, 8'h6E},
{8'h0B, 8'h26, 8'h60},
{8'h0B, 8'h1C, 8'h50},
{8'h0C, 8'h17, 8'h44},
{8'h0D, 8'h14, 8'h2F},
{8'h0C, 8'h13, 8'h30},
{8'h09, 8'h12, 8'h35},
{8'h07, 8'h11, 8'h3A},
{8'h01, 8'h0D, 8'h3A},
{8'h00, 8'h14, 8'h44},
{8'h01, 8'h1F, 8'h50},
{8'h06, 8'h27, 8'h5B},
{8'h11, 8'h38, 8'h88},
{8'h18, 8'h4B, 8'hA0},
{8'h1D, 8'h57, 8'hB0},
{8'h17, 8'h55, 8'hB4},
{8'h16, 8'h56, 8'hB8},
{8'h11, 8'h51, 8'hB5},
{8'h17, 8'h56, 8'hB8},
{8'h18, 8'h54, 8'hB6},
{8'h27, 8'h4B, 8'hA1},
{8'h21, 8'h41, 8'h8D},
{8'h16, 8'h2E, 8'h6D},
{8'h0D, 8'h1D, 8'h4F},
{8'h04, 8'h0E, 8'h3A},
{8'h04, 8'h08, 8'h36},
{8'h09, 8'h07, 8'h39},
{8'h10, 8'h0E, 8'h45},
{8'h07, 8'h19, 8'h5A},
{8'h0C, 8'h24, 8'h69},
{8'h19, 8'h34, 8'h76},
{8'h21, 8'h38, 8'h6E},
{8'hB1, 8'hBF, 8'hD5},
{8'hFF, 8'hFF, 8'hFF},
{8'hFE, 8'hF2, 8'hF3},
{8'hFF, 8'hF1, 8'hED},
{8'hFF, 8'hF9, 8'hF4},
{8'hFF, 8'hFD, 8'hF7},
{8'hFF, 8'hFD, 8'hF9},
{8'hFF, 8'hFE, 8'hFB},
{8'hFD, 8'hFB, 8'hFA},
{8'hF7, 8'hEF, 8'hF2},
{8'hDD, 8'hCC, 8'hD2},
{8'hE3, 8'hD3, 8'hDA},
{8'hFF, 8'hFD, 8'hFF},
{8'hFF, 8'hFF, 8'hFF},
{8'hFF, 8'hFE, 8'hFF},
{8'hFF, 8'hFD, 8'hFF},
{8'hFC, 8'hF8, 8'hFA},
{8'hFC, 8'hF8, 8'hF8},
{8'hFC, 8'hF8, 8'hF7},
{8'hFC, 8'hF8, 8'hF6},
{8'hFF, 8'hFB, 8'hFD},
{8'hFF, 8'hFE, 8'hFF},
{8'hFE, 8'hFE, 8'hFF},
{8'hFF, 8'hFC, 8'hFF},
{8'hFF, 8'hF8, 8'hFB},
{8'hF6, 8'hE6, 8'hE9},
{8'hEB, 8'hD5, 8'hDD},
{8'hB4, 8'hA3, 8'hB1},
{8'h07, 8'h08, 8'h1C},
{8'h05, 8'h03, 8'h17},
{8'h06, 8'h01, 8'h1B},
{8'h06, 8'h00, 8'h26},
{8'h02, 8'h04, 8'h22},
{8'h04, 8'h09, 8'h1A},
{8'h00, 8'h01, 8'h11},
{8'h04, 8'h04, 8'h1F},
{8'h24, 8'h16, 8'h2F},
{8'hA9, 8'h9D, 8'hA4},
{8'hFF, 8'hFD, 8'hF5},
{8'hFA, 8'hF7, 8'hED},
{8'hF8, 8'hF8, 8'hF4},
{8'hFD, 8'hFB, 8'hF6},
{8'hFD, 8'hF8, 8'hE1},
{8'hFE, 8'hF5, 8'hD1},
{8'hF9, 8'hEE, 8'hE0},
{8'hFC, 8'hF1, 8'hDF},
{8'hFA, 8'hE8, 8'hCD},
{8'hAA, 8'h7F, 8'h64},
{8'h6B, 8'h2E, 8'h1D},
{8'hD0, 8'hA3, 8'h8F},
{8'hFF, 8'hF8, 8'hE2},
{8'hF9, 8'hFD, 8'hE6},
{8'hF5, 8'hF3, 8'hDD},
{8'hA5, 8'hA2, 8'h85},
{8'hC6, 8'hC5, 8'hA0},
{8'hB5, 8'hB7, 8'h88},
{8'hDA, 8'hE1, 8'hAC},
{8'hEF, 8'hF8, 8'hC3},
{8'hEB, 8'hF3, 8'hC1},
{8'hF5, 8'hFE, 8'hD0},
{8'hC3, 8'hC4, 8'hB4},
{8'h7D, 8'h7D, 8'h73},
{8'h7F, 8'h7E, 8'h7B},
{8'h81, 8'h7F, 8'h83},
{8'h7F, 8'h7C, 8'h84},
{8'h7F, 8'h7C, 8'h84},
{8'h7F, 8'h7C, 8'h83},
{8'h7F, 8'h7C, 8'h83},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'h80, 8'h7C, 8'h7F},
{8'h8D, 8'h78, 8'h76},
{8'h9F, 8'h89, 8'h86},
{8'h96, 8'h82, 8'h7E},
{8'h94, 8'h81, 8'h7D},
{8'h9B, 8'h8B, 8'h86},
{8'hA8, 8'h9C, 8'h95},
{8'hB8, 8'hAD, 8'hA6},
{8'hB4, 8'hAD, 8'hA6},
{8'h92, 8'h8F, 8'h86},
{8'h7A, 8'h79, 8'h72},
{8'h79, 8'h7B, 8'h77},
{8'h7F, 8'h82, 8'h7D},
{8'h80, 8'h7E, 8'h76},
{8'h7E, 8'h73, 8'h64},
{8'h9F, 8'h89, 8'h70},
{8'hA7, 8'h8D, 8'h74},
{8'h51, 8'h56, 8'h6D},
{8'h2F, 8'h41, 8'h71},
{8'h2A, 8'h4F, 8'h96},
{8'h15, 8'h4D, 8'h9F},
{8'h05, 8'h4A, 8'h99},
{8'h03, 8'h4C, 8'h99},
{8'h09, 8'h49, 8'h99},
{8'h10, 8'h46, 8'h9B},
{8'h09, 8'h5A, 8'hB1},
{8'h0B, 8'h5F, 8'hB8},
{8'h0A, 8'h5C, 8'hBB},
{8'h0B, 8'h5A, 8'hBE},
{8'h0F, 8'h56, 8'hBE},
{8'h14, 8'h52, 8'hBB},
{8'h1A, 8'h4F, 8'hB8},
{8'h1C, 8'h4D, 8'hB6},
{8'h15, 8'h50, 8'hBD},
{8'h15, 8'h4F, 8'hBB},
{8'h17, 8'h4D, 8'hB6},
{8'h1B, 8'h4B, 8'hB1},
{8'h1E, 8'h48, 8'hAA},
{8'h1E, 8'h43, 8'hA1},
{8'h1E, 8'h3C, 8'h98},
{8'h1E, 8'h37, 8'h91},
{8'h15, 8'h39, 8'h8C},
{8'h0E, 8'h38, 8'h8C},
{8'h14, 8'h40, 8'h95},
{8'h19, 8'h4B, 8'hA1},
{8'h21, 8'h52, 8'hA6},
{8'h22, 8'h50, 8'hA0},
{8'h1A, 8'h42, 8'h8E},
{8'h16, 8'h3D, 8'h88},
{8'h12, 8'h41, 8'h97},
{8'h16, 8'h46, 8'hA1},
{8'h1B, 8'h47, 8'hA6},
{8'h1F, 8'h42, 8'hA1},
{8'h20, 8'h3B, 8'h92},
{8'h16, 8'h28, 8'h6F},
{8'h0E, 8'h1D, 8'h51},
{8'h00, 8'h08, 8'h30},
{8'h00, 8'h00, 8'h16},
{8'h00, 8'h00, 8'h1F},
{8'h00, 8'h00, 8'h21},
{8'h06, 8'h08, 8'h24},
{8'hC6, 8'hC2, 8'hC9},
{8'hF1, 8'hE0, 8'hDD},
{8'hF3, 8'hD2, 8'hD4},
{8'hF9, 8'hD2, 8'hDD},
{8'hEF, 8'hD9, 8'hDC},
{8'hEF, 8'hDE, 8'hDF},
{8'hF2, 8'hE3, 8'hE4},
{8'hF3, 8'hE8, 8'hE9},
{8'hEE, 8'hE1, 8'hE3},
{8'hE4, 8'hD0, 8'hD5},
{8'hD5, 8'hBC, 8'hC3},
{8'hEA, 8'hD0, 8'hD9},
{8'hFA, 8'hF1, 8'hF6},
{8'hF6, 8'hEA, 8'hF0},
{8'hEF, 8'hE3, 8'hE9},
{8'hEB, 8'hDD, 8'hE3},
{8'hE7, 8'hD6, 8'hDC},
{8'hE8, 8'hD5, 8'hDB},
{8'hE9, 8'hD5, 8'hDA},
{8'hE9, 8'hD5, 8'hD9},
{8'hF3, 8'hE0, 8'hE1},
{8'hF9, 8'hEF, 8'hF5},
{8'hFA, 8'hF4, 8'hFB},
{8'hF9, 8'hEB, 8'hF5},
{8'hF1, 8'hD9, 8'hDC},
{8'hED, 8'hD0, 8'hD3},
{8'hE8, 8'hD7, 8'hE5},
{8'h71, 8'h6E, 8'h89},
{8'h00, 8'h03, 8'h25},
{8'h04, 8'h03, 8'h16},
{8'h09, 8'h01, 8'h17},
{8'h07, 8'h00, 8'h29},
{8'h03, 8'h03, 8'h27},
{8'h07, 8'h0D, 8'h13},
{8'h45, 8'h43, 8'h3E},
{8'h16, 8'h04, 8'h0D},
{8'h24, 8'h0D, 8'h15},
{8'h99, 8'h83, 8'h78},
{8'hFF, 8'hF9, 8'hE2},
{8'hFD, 8'hF9, 8'hE7},
{8'hF9, 8'hFA, 8'hF7},
{8'hFB, 8'hF7, 8'hF3},
{8'hFF, 8'hF1, 8'hD7},
{8'hFB, 8'hDE, 8'hAF},
{8'hF0, 8'hD5, 8'hC1},
{8'hFD, 8'hF4, 8'hDE},
{8'hFF, 8'hF9, 8'hDF},
{8'h86, 8'h5E, 8'h4B},
{8'h49, 8'h04, 8'h00},
{8'h87, 8'h46, 8'h3A},
{8'hF8, 8'hE7, 8'hCF},
{8'hFA, 8'hFD, 8'hDD},
{8'hFC, 8'hF7, 8'hE6},
{8'hEA, 8'hE4, 8'hCD},
{8'hE1, 8'hDE, 8'hBA},
{8'hFA, 8'hFB, 8'hCD},
{8'hF4, 8'hF9, 8'hC6},
{8'hEC, 8'hF3, 8'hC2},
{8'hE9, 8'hF3, 8'hC5},
{8'hCF, 8'hD7, 8'hAF},
{8'h93, 8'h93, 8'h88},
{8'h7B, 8'h7A, 8'h75},
{8'h7C, 8'h7A, 8'h7A},
{8'h7F, 8'h7D, 8'h82},
{8'h7F, 8'h7C, 8'h84},
{8'h7F, 8'h7C, 8'h82},
{8'hFF, 8'hD7, 8'h00},
{8'h7F, 8'h7D, 8'h7E},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'h7F, 8'h7B, 8'h7E},
{8'h97, 8'h6E, 8'h6B},
{8'hCA, 8'hA1, 8'h9B},
{8'hF3, 8'hD4, 8'hCE},
{8'hF7, 8'hE3, 8'hDB},
{8'hFF, 8'hF0, 8'hE6},
{8'hFF, 8'hF6, 8'hEB},
{8'hFF, 8'hF8, 8'hEB},
{8'hFF, 8'hF7, 8'hEA},
{8'hFA, 8'hF0, 8'hE7},
{8'hD1, 8'hC8, 8'hC1},
{8'h93, 8'h87, 8'h83},
{8'h81, 8'h74, 8'h6D},
{8'h79, 8'h62, 8'h57},
{8'h4D, 8'h29, 8'h14},
{8'h91, 8'h5F, 8'h3D},
{8'hE6, 8'hAF, 8'h82},
{8'hE1, 8'hD3, 8'h90},
{8'h83, 8'h88, 8'h7D},
{8'h30, 8'h4C, 8'h91},
{8'h17, 8'h4E, 8'hC4},
{8'h0B, 8'h52, 8'hD0},
{8'h0B, 8'h54, 8'hB7},
{8'h19, 8'h5A, 8'h9B},
{8'h10, 8'h3F, 8'h71},
{8'h08, 8'h3A, 8'h8D},
{8'h16, 8'h53, 8'hAB},
{8'h11, 8'h53, 8'hAE},
{8'h13, 8'h5A, 8'hB5},
{8'h11, 8'h5B, 8'hB4},
{8'h12, 8'h5A, 8'hAE},
{8'h13, 8'h57, 8'hA6},
{8'h13, 8'h56, 8'hA4},
{8'h0E, 8'h59, 8'hB8},
{8'h0D, 8'h58, 8'hB6},
{8'h0F, 8'h57, 8'hB2},
{8'h12, 8'h56, 8'hAF},
{8'h18, 8'h59, 8'hB1},
{8'h1C, 8'h59, 8'hB1},
{8'h1D, 8'h57, 8'hB2},
{8'h1E, 8'h57, 8'hB2},
{8'h1C, 8'h57, 8'hAF},
{8'h22, 8'h5B, 8'hB0},
{8'h22, 8'h56, 8'hA6},
{8'h1F, 8'h4B, 8'h92},
{8'h15, 8'h31, 8'h6B},
{8'h00, 8'h0E, 8'h3A},
{8'h00, 8'h00, 8'h1D},
{8'h00, 8'h00, 8'h17},
{8'h00, 8'h00, 8'h26},
{8'h00, 8'h00, 8'h22},
{8'h00, 8'h02, 8'h18},
{8'h00, 8'h03, 8'h0F},
{8'h03, 8'h0B, 8'h0F},
{8'h0F, 8'h15, 8'h17},
{8'h1A, 8'h1F, 8'h25},
{8'h1B, 8'h1C, 8'h26},
{8'h29, 8'h26, 8'h1C},
{8'h36, 8'h32, 8'h30},
{8'h4B, 8'h48, 8'h53},
{8'h84, 8'h7F, 8'h84},
{8'hBD, 8'hB6, 8'hAA},
{8'hED, 8'hDB, 8'hCC},
{8'hEB, 8'hCC, 8'hCF},
{8'hEF, 8'hC6, 8'hDD},
{8'hE6, 8'hC9, 8'hD5},
{8'hE6, 8'hCC, 8'hD5},
{8'hE7, 8'hCF, 8'hD7},
{8'hE8, 8'hD3, 8'hD8},
{8'hE7, 8'hD0, 8'hD6},
{8'hE1, 8'hC7, 8'hCD},
{8'hD8, 8'hB8, 8'hBE},
{8'hE5, 8'hC3, 8'hCA},
{8'hE6, 8'hD1, 8'hD4},
{8'hE4, 8'hD0, 8'hD2},
{8'hE3, 8'hCC, 8'hD2},
{8'hE5, 8'hCB, 8'hD1},
{8'hE8, 8'hCC, 8'hD4},
{8'hEA, 8'hCB, 8'hD5},
{8'hEB, 8'hCA, 8'hD6},
{8'hEB, 8'hC9, 8'hD4},
{8'hE8, 8'hC5, 8'hC6},
{8'hE6, 8'hD0, 8'hD9},
{8'hE2, 8'hD4, 8'hE6},
{8'hE3, 8'hCE, 8'hDC},
{8'hEF, 8'hCD, 8'hD0},
{8'hEC, 8'hCB, 8'hCE},
{8'hD0, 8'hC4, 8'hD3},
{8'h30, 8'h39, 8'h59},
{8'h04, 8'h0F, 8'h39},
{8'h04, 8'h03, 8'h15},
{8'h0C, 8'h01, 8'h14},
{8'h09, 8'h00, 8'h2C},
{8'h01, 8'h00, 8'h29},
{8'h07, 8'h0D, 8'h0D},
{8'hB5, 8'hAC, 8'h99},
{8'hA1, 8'h86, 8'h86},
{8'hB3, 8'hA9, 8'hAB},
{8'hF4, 8'hEA, 8'hD3},
{8'hFF, 8'hEC, 8'hBE},
{8'hFE, 8'hE9, 8'hBF},
{8'hF8, 8'hEA, 8'hD6},
{8'hFA, 8'hEE, 8'hE4},
{8'hF8, 8'hE1, 8'hC5},
{8'hF0, 8'hC0, 8'h91},
{8'hEE, 8'hCB, 8'hB1},
{8'hFF, 8'hF2, 8'hD8},
{8'hFF, 8'hFB, 8'hE4},
{8'h8E, 8'h69, 8'h5F},
{8'h45, 8'h03, 8'h01},
{8'h79, 8'h30, 8'h29},
{8'hC4, 8'h9F, 8'h83},
{8'hFF, 8'hFF, 8'hD6},
{8'hFD, 8'hF6, 8'hE7},
{8'hFE, 8'hF5, 8'hE0},
{8'hDE, 8'hD9, 8'hB7},
{8'hEB, 8'hEC, 8'hC0},
{8'hEE, 8'hF3, 8'hC1},
{8'hEB, 8'hF2, 8'hC4},
{8'hE9, 8'hF0, 8'hCA},
{8'h92, 8'h9A, 8'h7C},
{8'h7D, 8'h7D, 8'h78},
{8'h7F, 8'h7D, 8'h7D},
{8'h80, 8'h7E, 8'h81},
{8'h7D, 8'h7B, 8'h81},
{8'h7F, 8'h7D, 8'h82},
{8'hFF, 8'hD7, 8'h00},
{8'h7F, 8'h7E, 8'h7A},
{8'h7F, 8'h7E, 8'h78},
{8'h80, 8'h7E, 8'h82},
{8'h7F, 8'h7D, 8'h81},
{8'h7F, 8'h7C, 8'h81},
{8'h80, 8'h7D, 8'h81},
{8'h7F, 8'h7C, 8'h80},
{8'h80, 8'h7C, 8'h80},
{8'h81, 8'h7C, 8'h80},
{8'h82, 8'h7C, 8'h7F},
{8'h90, 8'h6F, 8'h6F},
{8'h95, 8'h73, 8'h71},
{8'hA8, 8'h8C, 8'h88},
{8'hBC, 8'hA7, 8'hA0},
{8'hC5, 8'hB0, 8'hA7},
{8'hE0, 8'hCF, 8'hC3},
{8'hFF, 8'hF7, 8'hEA},
{8'hFF, 8'hF2, 8'hE4},
{8'hFF, 8'hF0, 8'hEA},
{8'hFF, 8'hF2, 8'hEF},
{8'hF8, 8'hE7, 8'hE4},
{8'hD8, 8'hC4, 8'hBE},
{8'hD7, 8'hBD, 8'hB1},
{8'hDA, 8'hC2, 8'hAC},
{8'hC7, 8'h97, 8'h77},
{8'h97, 8'h5A, 8'h30},
{8'hCB, 8'h96, 8'h37},
{8'hFA, 8'hE2, 8'h88},
{8'h94, 8'h9C, 8'h80},
{8'h2C, 8'h51, 8'h9B},
{8'h1B, 8'h56, 8'hBE},
{8'h17, 8'h52, 8'hC7},
{8'h1D, 8'h4C, 8'hB9},
{8'h26, 8'h4B, 8'h9B},
{8'h0B, 8'h1E, 8'h69},
{8'h1D, 8'h3A, 8'h8C},
{8'h26, 8'h53, 8'hAE},
{8'h18, 8'h50, 8'hB5},
{8'h12, 8'h53, 8'hBF},
{8'h10, 8'h54, 8'hC2},
{8'h12, 8'h54, 8'hC4},
{8'h13, 8'h56, 8'hC1},
{8'h15, 8'h58, 8'hAB},
{8'h17, 8'h59, 8'hAC},
{8'h14, 8'h55, 8'hAF},
{8'h15, 8'h54, 8'hB4},
{8'h16, 8'h53, 8'hB8},
{8'h18, 8'h52, 8'hBB},
{8'h18, 8'h52, 8'hBD},
{8'h18, 8'h50, 8'hBA},
{8'h19, 8'h45, 8'h96},
{8'h0A, 8'h34, 8'h7B},
{8'h00, 8'h1B, 8'h55},
{8'h05, 8'h13, 8'h3F},
{8'h23, 8'h26, 8'h45},
{8'h39, 8'h39, 8'h47},
{8'h54, 8'h4F, 8'h4F},
{8'h76, 8'h6B, 8'h61},
{8'h84, 8'h80, 8'h71},
{8'hA0, 8'h9E, 8'h91},
{8'hB5, 8'hB3, 8'hAD},
{8'hB3, 8'hB5, 8'hB2},
{8'h99, 8'hA0, 8'h96},
{8'hB2, 8'hBD, 8'hA4},
{8'hAC, 8'hBC, 8'h95},
{8'hA7, 8'hB8, 8'h89},
{8'hC0, 8'hC0, 8'h92},
{8'hD8, 8'hD5, 8'hB9},
{8'hE6, 8'hE1, 8'hD7},
{8'hF4, 8'hED, 8'hE6},
{8'hC3, 8'hB9, 8'hAC},
{8'hE1, 8'hD0, 8'hC6},
{8'hE6, 8'hC9, 8'hD2},
{8'hEC, 8'hC9, 8'hE2},
{8'hE9, 8'hCB, 8'hD9},
{8'hEA, 8'hCE, 8'hD9},
{8'hE8, 8'hCD, 8'hD7},
{8'hE5, 8'hCB, 8'hD3},
{8'hE5, 8'hCB, 8'hD2},
{8'hEB, 8'hCD, 8'hD4},
{8'hE9, 8'hC8, 8'hCF},
{8'hEE, 8'hCB, 8'hD3},
{8'hE7, 8'hCC, 8'hCD},
{8'hE7, 8'hCC, 8'hCF},
{8'hE7, 8'hCB, 8'hD0},
{8'hE8, 8'hCB, 8'hD3},
{8'hE9, 8'hCB, 8'hD5},
{8'hEB, 8'hCA, 8'hD7},
{8'hEC, 8'hC9, 8'hD8},
{8'hED, 8'hCA, 8'hD7},
{8'hE8, 8'hCE, 8'hD3},
{8'hE1, 8'hCC, 8'hDA},
{8'hE0, 8'hC9, 8'hDE},
{8'hE6, 8'hC6, 8'hD2},
{8'hEE, 8'hC9, 8'hC9},
{8'hE9, 8'hD0, 8'hD3},
{8'h8C, 8'h8F, 8'hA9},
{8'h24, 8'h3E, 8'h70},
{8'h10, 8'h1A, 8'h4B},
{8'h03, 8'h02, 8'h18},
{8'h09, 8'h04, 8'h15},
{8'h06, 8'h01, 8'h27},
{8'h01, 8'h00, 8'h21},
{8'h4F, 8'h50, 8'h4E},
{8'hEA, 8'hE6, 8'hC9},
{8'hFF, 8'hFC, 8'hDE},
{8'hFF, 8'hF9, 8'hE3},
{8'hFD, 8'hE0, 8'hBD},
{8'hF2, 8'hC4, 8'h94},
{8'hD8, 8'hAA, 8'h7F},
{8'hEB, 8'hCF, 8'hB5},
{8'hFD, 8'hF5, 8'hE4},
{8'hEB, 8'hC2, 8'hAA},
{8'h9A, 8'h59, 8'h36},
{8'hBF, 8'h98, 8'h7F},
{8'hFF, 8'hFC, 8'hE1},
{8'hFF, 8'hFD, 8'hE5},
{8'hA7, 8'h84, 8'h78},
{8'h46, 8'h02, 8'h03},
{8'h7C, 8'h31, 8'h29},
{8'hCC, 8'hA6, 8'h88},
{8'hF2, 8'hEE, 8'hC2},
{8'hFD, 8'hF9, 8'hE8},
{8'hF6, 8'hEF, 8'hDC},
{8'hF8, 8'hF4, 8'hDB},
{8'hD7, 8'hD2, 8'hB2},
{8'hED, 8'hEC, 8'hC6},
{8'hEE, 8'hF2, 8'hCB},
{8'hEE, 8'hF8, 8'hD0},
{8'hCA, 8'hD7, 8'hB2},
{8'h7E, 8'h7D, 8'h78},
{8'h78, 8'h76, 8'h79},
{8'h82, 8'h80, 8'h86},
{8'h80, 8'h7D, 8'h85},
{8'h7F, 8'h7D, 8'h7F},
{8'h7F, 8'h7E, 8'h7C},
{8'h7F, 8'h7E, 8'h7B},
{8'h7F, 8'h7E, 8'h7B},
{8'h7D, 8'h7C, 8'h83},
{8'h7E, 8'h7E, 8'h84},
{8'h80, 8'h7E, 8'h84},
{8'h80, 8'h7C, 8'h82},
{8'h7E, 8'h79, 8'h7D},
{8'h80, 8'h7A, 8'h7E},
{8'h83, 8'h7D, 8'h7E},
{8'h84, 8'h7D, 8'h80},
{8'h7F, 8'h7D, 8'h84},
{8'h7F, 8'h7F, 8'h85},
{8'h77, 8'h78, 8'h79},
{8'h71, 8'h6F, 8'h6B},
{8'h74, 8'h6E, 8'h67},
{8'h9D, 8'h8F, 8'h86},
{8'hE7, 8'hD5, 8'hCB},
{8'hFF, 8'hEB, 8'hE0},
{8'hFF, 8'hEF, 8'hE8},
{8'hFD, 8'hF0, 8'hEA},
{8'hFD, 8'hF3, 8'hED},
{8'hFF, 8'hF6, 8'hF0},
{8'hFF, 8'hF8, 8'hEF},
{8'hFF, 8'hF4, 8'hE8},
{8'hFF, 8'hF9, 8'hE9},
{8'hDD, 8'hC4, 8'hB1},
{8'hA0, 8'h44, 8'h3B},
{8'hCE, 8'h8E, 8'h49},
{8'hFB, 8'hE7, 8'h70},
{8'h7C, 8'h86, 8'h93},
{8'h1F, 8'h51, 8'h98},
{8'h10, 8'h54, 8'hC5},
{8'h10, 8'h53, 8'hC3},
{8'h1B, 8'h58, 8'h9D},
{8'h11, 8'h20, 8'h60},
{8'h0B, 8'h21, 8'h69},
{8'h1F, 8'h53, 8'hA6},
{8'h14, 8'h56, 8'hB3},
{8'h0B, 8'h57, 8'hBB},
{8'h09, 8'h57, 8'hBC},
{8'h0A, 8'h56, 8'hB9},
{8'h0C, 8'h55, 8'hB4},
{8'h0D, 8'h58, 8'hAC},
{8'h11, 8'h57, 8'hAF},
{8'h19, 8'h56, 8'hB4},
{8'h20, 8'h51, 8'hB3},
{8'h21, 8'h46, 8'hA2},
{8'h1D, 8'h39, 8'h89},
{8'h11, 8'h21, 8'h63},
{8'h03, 8'h10, 8'h47},
{8'h03, 8'h00, 8'h20},
{8'h1F, 8'h1A, 8'h2C},
{8'h65, 8'h63, 8'h66},
{8'hC5, 8'hC3, 8'hC3},
{8'hE9, 8'hE8, 8'hEB},
{8'hF2, 8'hF3, 8'hF4},
{8'hFA, 8'hFD, 8'hF3},
{8'hFA, 8'hFF, 8'hEA},
{8'hFF, 8'hFD, 8'hEF},
{8'hFE, 8'hF9, 8'hF0},
{8'hFF, 8'hFC, 8'hFA},
{8'hFE, 8'hFA, 8'hF8},
{8'hF2, 8'hF3, 8'hE9},
{8'hE5, 8'hEA, 8'hD0},
{8'hB9, 8'hC2, 8'h95},
{8'hDB, 8'hE7, 8'hAF},
{8'hC5, 8'hD0, 8'h9B},
{8'hC2, 8'hC9, 8'h9D},
{8'hAD, 8'hAD, 8'h90},
{8'hED, 8'hE5, 8'hD8},
{8'hC7, 8'hB6, 8'hB8},
{8'hE2, 8'hCA, 8'hD4},
{8'hE9, 8'hCC, 8'hD8},
{8'hE8, 8'hCA, 8'hD4},
{8'hE5, 8'hCC, 8'hD5},
{8'hE7, 8'hCD, 8'hD6},
{8'hE7, 8'hCD, 8'hD6},
{8'hE7, 8'hCC, 8'hD5},
{8'hE7, 8'hCC, 8'hD5},
{8'hE7, 8'hCA, 8'hD4},
{8'hE7, 8'hC9, 8'hD3},
{8'hE7, 8'hC8, 8'hD3},
{8'hEA, 8'hCA, 8'hD0},
{8'hEA, 8'hCB, 8'hD1},
{8'hE9, 8'hCC, 8'hD5},
{8'hE7, 8'hCD, 8'hD7},
{8'hE5, 8'hCB, 8'hD6},
{8'hE5, 8'hCB, 8'hD6},
{8'hE6, 8'hCA, 8'hD5},
{8'hE6, 8'hCB, 8'hD4},
{8'hD5, 8'hD0, 8'hD9},
{8'hDF, 8'hCB, 8'hDE},
{8'hEF, 8'hC7, 8'hDB},
{8'hF5, 8'hC7, 8'hCE},
{8'hE9, 8'hCD, 8'hC9},
{8'hC7, 8'hCC, 8'hD9},
{8'h36, 8'h5C, 8'h94},
{8'h1A, 8'h4E, 8'hA8},
{8'h14, 8'h16, 8'h4C},
{8'h00, 8'h00, 8'h21},
{8'h00, 8'h05, 8'h18},
{8'h00, 8'h05, 8'h14},
{8'h0D, 8'h0E, 8'h1E},
{8'hDC, 8'hD6, 8'hD4},
{8'hFF, 8'hF8, 8'hCE},
{8'hEF, 8'hE3, 8'h93},
{8'hDF, 8'hC1, 8'h7C},
{8'hE9, 8'hB9, 8'h89},
{8'hD0, 8'h9C, 8'h84},
{8'h9B, 8'h71, 8'h65},
{8'hF4, 8'hE3, 8'hD6},
{8'hFF, 8'hF5, 8'hE2},
{8'hD9, 8'hA0, 8'h8C},
{8'h79, 8'h20, 8'h0D},
{8'hB0, 8'h87, 8'h78},
{8'hFF, 8'hFC, 8'hE4},
{8'hFF, 8'hFD, 8'hE0},
{8'hBB, 8'h9A, 8'h80},
{8'h53, 8'h0F, 8'h02},
{8'h75, 8'h31, 8'h1D},
{8'hF2, 8'hDC, 8'hB8},
{8'hD8, 8'hDF, 8'hB1},
{8'hF4, 8'hF7, 8'hDB},
{8'hFA, 8'hF8, 8'hE6},
{8'hFB, 8'hEF, 8'hE5},
{8'hF5, 8'hE5, 8'hDE},
{8'hD2, 8'hC2, 8'hB3},
{8'hF0, 8'hEC, 8'hCD},
{8'hF1, 8'hFB, 8'hC9},
{8'hE0, 8'hF1, 8'hB5},
{8'h82, 8'h84, 8'h73},
{8'h7D, 8'h7C, 8'h7B},
{8'h7E, 8'h7B, 8'h85},
{8'h7D, 8'h7A, 8'h82},
{8'h7E, 8'h7D, 8'h7C},
{8'h7F, 8'h7E, 8'h79},
{8'hFF, 8'hD7, 8'h00},
{8'h7F, 8'h7C, 8'h88},
{8'h7B, 8'h7D, 8'h7E},
{8'h7F, 8'h81, 8'h83},
{8'h81, 8'h82, 8'h82},
{8'h7E, 8'h7F, 8'h7E},
{8'h7E, 8'h7E, 8'h7C},
{8'h7F, 8'h7D, 8'h7A},
{8'h7E, 8'h7C, 8'h78},
{8'h7F, 8'h7A, 8'h77},
{8'h82, 8'h78, 8'h7B},
{8'h81, 8'h75, 8'h78},
{8'h86, 8'h7C, 8'h7A},
{8'hAD, 8'hA4, 8'h9F},
{8'hE3, 8'hDA, 8'hD1},
{8'hF4, 8'hE5, 8'hDA},
{8'hF1, 8'hD9, 8'hCE},
{8'hFF, 8'hE9, 8'hDD},
{8'hFF, 8'hF1, 8'hDE},
{8'hFB, 8'hE7, 8'hD6},
{8'hF7, 8'hE6, 8'hD9},
{8'hFA, 8'hEE, 8'hE5},
{8'hF8, 8'hEF, 8'hE6},
{8'hFC, 8'hF2, 8'hEA},
{8'hFC, 8'hF2, 8'hE9},
{8'hFF, 8'hF8, 8'hE8},
{8'hCA, 8'h94, 8'h78},
{8'h92, 8'h45, 8'h2E},
{8'hEC, 8'hBF, 8'h4A},
{8'hD8, 8'hCF, 8'h8C},
{8'h2D, 8'h4E, 8'h94},
{8'h0B, 8'h53, 8'hB7},
{8'h0C, 8'h5C, 8'hB6},
{8'h18, 8'h56, 8'hB5},
{8'h15, 8'h1C, 8'h4D},
{8'h03, 8'h0B, 8'h3F},
{8'h1D, 8'h3A, 8'h7B},
{8'h23, 8'h4A, 8'h97},
{8'h20, 8'h4D, 8'hA4},
{8'h20, 8'h4C, 8'hA7},
{8'h21, 8'h4A, 8'hA6},
{8'h23, 8'h49, 8'hA4},
{8'h1F, 8'h45, 8'hA5},
{8'h19, 8'h3D, 8'h96},
{8'h11, 8'h2E, 8'h7A},
{8'h09, 8'h1F, 8'h59},
{8'h00, 8'h0A, 8'h2F},
{8'h00, 8'h06, 8'h16},
{8'h14, 8'h1D, 8'h1A},
{8'h51, 8'h5C, 8'h51},
{8'hA1, 8'hA6, 8'h9C},
{8'hD4, 8'hDA, 8'hC6},
{8'hF7, 8'hFC, 8'hE3},
{8'hFF, 8'hFF, 8'hF3},
{8'hFF, 8'hFF, 8'hFA},
{8'hFD, 8'hFB, 8'hFE},
{8'hF7, 8'hF5, 8'hF3},
{8'hF4, 8'hF1, 8'hE7},
{8'hF5, 8'hF4, 8'hDA},
{8'hE7, 8'hE5, 8'hD1},
{8'hFA, 8'hF6, 8'hEC},
{8'hF9, 8'hF6, 8'hF3},
{8'hF8, 8'hF8, 8'hF1},
{8'hF6, 8'hF9, 8'hE7},
{8'hB6, 8'hBD, 8'h9C},
{8'hC8, 8'hD1, 8'hA7},
{8'hC7, 8'hCF, 8'hA0},
{8'hAD, 8'hB2, 8'h8B},
{8'h9A, 8'h9A, 8'h7D},
{8'hF0, 8'hE9, 8'hD8},
{8'hD1, 8'hC3, 8'hBC},
{8'hD8, 8'hC4, 8'hC1},
{8'hE7, 8'hCF, 8'hCE},
{8'hE6, 8'hCC, 8'hCB},
{8'hE5, 8'hCB, 8'hD3},
{8'hE9, 8'hCE, 8'hD7},
{8'hE8, 8'hCE, 8'hD7},
{8'hE4, 8'hCB, 8'hD4},
{8'hE5, 8'hCC, 8'hD5},
{8'hE5, 8'hCE, 8'hD6},
{8'hE1, 8'hCA, 8'hD2},
{8'hDC, 8'hC6, 8'hCD},
{8'hEA, 8'hCC, 8'hD4},
{8'hEC, 8'hCE, 8'hD6},
{8'hEC, 8'hCF, 8'hD7},
{8'hEB, 8'hCF, 8'hD8},
{8'hE7, 8'hCB, 8'hD2},
{8'hE7, 8'hCB, 8'hD2},
{8'hE8, 8'hCB, 8'hD0},
{8'hE9, 8'hCB, 8'hCE},
{8'hF2, 8'hCC, 8'hC3},
{8'hF6, 8'hCB, 8'hCF},
{8'hF0, 8'hC4, 8'hD5},
{8'hEE, 8'hCC, 8'hDE},
{8'hD7, 8'hCE, 8'hE1},
{8'h65, 8'h7D, 8'hA1},
{8'h1C, 8'h50, 8'h99},
{8'h12, 8'h50, 8'hB2},
{8'h0D, 8'h11, 8'h43},
{8'h00, 8'h01, 8'h21},
{8'h00, 8'h04, 8'h17},
{8'h00, 8'h05, 8'h15},
{8'h0E, 8'h10, 8'h1D},
{8'hB8, 8'hB1, 8'hAB},
{8'hE3, 8'hD4, 8'hAA},
{8'hD2, 8'hBF, 8'h78},
{8'hDE, 8'hD1, 8'h92},
{8'hF3, 8'hDC, 8'hAC},
{8'hFB, 8'hE2, 8'hC5},
{8'hEB, 8'hD8, 8'hC5},
{8'hFB, 8'hF3, 8'hE2},
{8'hF8, 8'hF1, 8'hDB},
{8'hCE, 8'hAC, 8'h94},
{8'hAB, 8'h75, 8'h5F},
{8'hBF, 8'h9C, 8'h8D},
{8'hFE, 8'hF4, 8'hDF},
{8'hFF, 8'hFF, 8'hE5},
{8'hCF, 8'hB9, 8'h9F},
{8'h5E, 8'h28, 8'h12},
{8'h8E, 8'h5A, 8'h42},
{8'hFC, 8'hEE, 8'hC3},
{8'hE7, 8'hF3, 8'hBD},
{8'hDC, 8'hD5, 8'hB8},
{8'hF6, 8'hEA, 8'hD5},
{8'hFF, 8'hEE, 8'hE1},
{8'hFD, 8'hE5, 8'hDA},
{8'hE5, 8'hD0, 8'hBF},
{8'hDB, 8'hCC, 8'hAD},
{8'hF7, 8'hF3, 8'hC4},
{8'hE2, 8'hE6, 8'hAE},
{8'h82, 8'h84, 8'h70},
{8'h7E, 8'h7D, 8'h79},
{8'h80, 8'h7C, 8'h86},
{8'h7D, 8'h7A, 8'h83},
{8'h7F, 8'h7D, 8'h7E},
{8'h7F, 8'h7E, 8'h7A},
{8'hFF, 8'hD7, 8'h00},
{8'h7F, 8'h7C, 8'h87},
{8'h82, 8'h80, 8'h7D},
{8'h80, 8'h7E, 8'h7A},
{8'h7D, 8'h79, 8'h74},
{8'h7C, 8'h78, 8'h73},
{8'h8A, 8'h85, 8'h7E},
{8'h91, 8'h8B, 8'h83},
{8'h99, 8'h91, 8'h89},
{8'h9D, 8'h94, 8'h8D},
{8'hA6, 8'h91, 8'h90},
{8'hC6, 8'hB4, 8'hB2},
{8'hF1, 8'hE3, 8'hDE},
{8'hFF, 8'hF6, 8'hEE},
{8'hFF, 8'hF5, 8'hE9},
{8'hFF, 8'hEC, 8'hDF},
{8'hFF, 8'hE8, 8'hDA},
{8'hF1, 8'hD4, 8'hC6},
{8'hDE, 8'hC4, 8'hAE},
{8'hEF, 8'hD8, 8'hC3},
{8'hFB, 8'hEC, 8'hDB},
{8'hFC, 8'hF4, 8'hE8},
{8'hFE, 8'hF6, 8'hEC},
{8'hFB, 8'hF2, 8'hE8},
{8'hFB, 8'hEF, 8'hE6},
{8'hFE, 8'hFA, 8'hEB},
{8'hE6, 8'hC5, 8'hA6},
{8'h93, 8'h3D, 8'h39},
{8'hD2, 8'h8D, 8'h2B},
{8'hF0, 8'hDA, 8'h6E},
{8'h34, 8'h52, 8'h86},
{8'h08, 8'h58, 8'hB1},
{8'h0B, 8'h59, 8'hC2},
{8'h16, 8'h48, 8'hAD},
{8'h10, 8'h0F, 8'h30},
{8'h04, 8'h03, 8'h25},
{8'h03, 8'h06, 8'h33},
{8'h05, 8'h0C, 8'h41},
{8'h07, 8'h0E, 8'h48},
{8'h06, 8'h0C, 8'h48},
{8'h05, 8'h08, 8'h44},
{8'h01, 8'h04, 8'h3D},
{8'h00, 8'h04, 8'h35},
{8'h00, 8'h00, 8'h26},
{8'h00, 8'h04, 8'h18},
{8'h26, 8'h28, 8'h29},
{8'h54, 8'h5A, 8'h4B},
{8'h94, 8'h99, 8'h82},
{8'hD1, 8'hD6, 8'hBB},
{8'hFF, 8'hFF, 8'hE5},
{8'hF4, 8'hFE, 8'hD5},
{8'hE6, 8'hF3, 8'hC0},
{8'hE2, 8'hED, 8'hBC},
{8'hF6, 8'hFA, 8'hDA},
{8'hF9, 8'hF9, 8'hED},
{8'hF7, 8'hF3, 8'hF4},
{8'hF4, 8'hED, 8'hED},
{8'hEF, 8'hE8, 8'hDE},
{8'hDF, 8'hE1, 8'hB7},
{8'hE3, 8'hE4, 8'hC1},
{8'hFB, 8'hFA, 8'hE6},
{8'hF9, 8'hF7, 8'hF0},
{8'hF3, 8'hF2, 8'hED},
{8'hF7, 8'hF8, 8'hF0},
{8'hEE, 8'hF0, 8'hDF},
{8'hC4, 8'hC8, 8'hB0},
{8'hC6, 8'hC9, 8'hA9},
{8'hB1, 8'hB2, 8'h95},
{8'hDC, 8'hD9, 8'hC3},
{8'hF3, 8'hEC, 8'hDC},
{8'hE6, 8'hDB, 8'hD1},
{8'hC9, 8'hBA, 8'hB2},
{8'hE1, 8'hCF, 8'hC8},
{8'hE7, 8'hD3, 8'hCD},
{8'hE7, 8'hCB, 8'hD4},
{8'hEA, 8'hCF, 8'hD8},
{8'hE7, 8'hCE, 8'hD6},
{8'hE2, 8'hCC, 8'hD3},
{8'hE7, 8'hD5, 8'hDC},
{8'hE9, 8'hDA, 8'hDF},
{8'hE1, 8'hD5, 8'hD9},
{8'hD5, 8'hC9, 8'hCD},
{8'hE2, 8'hC8, 8'hD3},
{8'hE5, 8'hCA, 8'hD5},
{8'hE7, 8'hCB, 8'hD4},
{8'hE7, 8'hCB, 8'hD2},
{8'hE6, 8'hCB, 8'hD0},
{8'hE7, 8'hCD, 8'hD2},
{8'hE9, 8'hD0, 8'hD4},
{8'hEB, 8'hD0, 8'hD3},
{8'hFE, 8'hCA, 8'hC1},
{8'hFA, 8'hCD, 8'hD2},
{8'hEB, 8'hCE, 8'hE9},
{8'hBC, 8'hB8, 8'hE1},
{8'h60, 8'h75, 8'hAA},
{8'h20, 8'h4D, 8'h90},
{8'h19, 8'h58, 8'hB1},
{8'h0E, 8'h4E, 8'hB3},
{8'h06, 8'h0B, 8'h38},
{8'h01, 8'h03, 8'h22},
{8'h00, 8'h04, 8'h17},
{8'h00, 8'h04, 8'h11},
{8'h10, 8'h10, 8'h16},
{8'hC4, 8'hBD, 8'hB1},
{8'hF6, 8'hE9, 8'hC2},
{8'hE3, 8'hD4, 8'h98},
{8'hD5, 8'hD7, 8'hA1},
{8'hE5, 8'hE2, 8'hB7},
{8'hF6, 8'hF0, 8'hD2},
{8'hE4, 8'hE1, 8'hCC},
{8'hFD, 8'hFD, 8'hEC},
{8'hF3, 8'hF3, 8'hDE},
{8'hE0, 8'hD6, 8'hBF},
{8'hFF, 8'hFC, 8'hE6},
{8'hE9, 8'hD8, 8'hCD},
{8'hF9, 8'hF3, 8'hE2},
{8'hFD, 8'hFA, 8'hE2},
{8'hDD, 8'hCD, 8'hB2},
{8'hA6, 8'h84, 8'h68},
{8'hC1, 8'hA3, 8'h80},
{8'hFA, 8'hF7, 8'hC3},
{8'hE5, 8'hFA, 8'hBD},
{8'hEF, 8'hE6, 8'hC2},
{8'hE0, 8'hD0, 8'hB3},
{8'hEA, 8'hD2, 8'hBB},
{8'hFA, 8'hE2, 8'hCD},
{8'hF2, 8'hDD, 8'hC4},
{8'hC3, 8'hAF, 8'h8C},
{8'hF7, 8'hED, 8'hBE},
{8'hF4, 8'hF0, 8'hBB},
{8'hB4, 8'hB6, 8'h9D},
{8'h81, 8'h80, 8'h79},
{8'h7E, 8'h7B, 8'h83},
{8'h79, 8'h76, 8'h80},
{8'hFF, 8'hD7, 8'h00},
{8'h7F, 8'h7E, 8'h7B},
{8'hFF, 8'hD7, 8'h00},
{8'h7F, 8'h7C, 8'h85},
{8'h85, 8'h75, 8'h72},
{8'h8F, 8'h7F, 8'h7C},
{8'hC2, 8'hB2, 8'hAE},
{8'hE7, 8'hD8, 8'hD2},
{8'hF2, 8'hE6, 8'hE0},
{8'hF4, 8'hE4, 8'hDD},
{8'hF6, 8'hE3, 8'hDB},
{8'hF8, 8'hE4, 8'hDD},
{8'hF6, 8'hDA, 8'hD6},
{8'hFE, 8'hE6, 8'hE0},
{8'hFF, 8'hF5, 8'hEC},
{8'hFA, 8'hE2, 8'hD7},
{8'hE2, 8'hC7, 8'hBA},
{8'hDB, 8'hBC, 8'hAD},
{8'hDA, 8'hB2, 8'hA4},
{8'hE2, 8'hBA, 8'hAA},
{8'hF4, 8'hE5, 8'hD6},
{8'hFD, 8'hF2, 8'hE4},
{8'hFF, 8'hF5, 8'hE9},
{8'hFC, 8'hF0, 8'hE5},
{8'hFC, 8'hF0, 8'hE3},
{8'hFF, 8'hF2, 8'hE2},
{8'hFF, 8'hED, 8'hD9},
{8'hF8, 8'hDE, 8'hC7},
{8'hD8, 8'hA5, 8'h8A},
{8'h9D, 8'h43, 8'h40},
{8'hD6, 8'h87, 8'h46},
{8'hDB, 8'hC6, 8'h6C},
{8'h28, 8'h54, 8'h88},
{8'h07, 8'h5D, 8'hB7},
{8'h14, 8'h4E, 8'hCB},
{8'h1E, 8'h33, 8'h84},
{8'h05, 8'h02, 8'h1E},
{8'h08, 8'h03, 8'h22},
{8'h04, 8'h03, 8'h20},
{8'h00, 8'h00, 8'h19},
{8'h00, 8'h00, 8'h11},
{8'h00, 8'h00, 8'h0E},
{8'h16, 8'h15, 8'h1C},
{8'h3A, 8'h3A, 8'h3A},
{8'h5B, 8'h61, 8'h4D},
{8'h97, 8'h9E, 8'h82},
{8'hBC, 8'hC5, 8'h9E},
{8'hDD, 8'hE6, 8'hBB},
{8'hED, 8'hF4, 8'hCC},
{8'hF4, 8'hF7, 8'hDC},
{8'hF8, 8'hF7, 8'hED},
{8'hF5, 8'hF3, 8'hF0},
{8'hE6, 8'hEF, 8'hCD},
{8'hDF, 8'hEC, 8'hBF},
{8'hE3, 8'hEC, 8'hC2},
{8'hDF, 8'hE3, 8'hC6},
{8'hE7, 8'hE6, 8'hDB},
{8'hEC, 8'hE6, 8'hE3},
{8'hEF, 8'hE7, 8'hDF},
{8'hE7, 8'hE0, 8'hCB},
{8'hE5, 8'hEB, 8'hB4},
{8'hEB, 8'hF0, 8'hC2},
{8'hF2, 8'hF4, 8'hD9},
{8'hFC, 8'hFC, 8'hF1},
{8'hF7, 8'hF6, 8'hF3},
{8'hF6, 8'hF5, 8'hF3},
{8'hFB, 8'hFA, 8'hF3},
{8'hEB, 8'hEB, 8'hDE},
{8'hC4, 8'hC1, 8'hB1},
{8'hE4, 8'hE1, 8'hD1},
{8'hF6, 8'hF0, 8'hE4},
{8'hF0, 8'hE8, 8'hDF},
{8'hF1, 8'hE7, 8'hE3},
{8'hC8, 8'hBB, 8'hBB},
{8'hDA, 8'hCC, 8'hCD},
{8'hEB, 8'hDB, 8'hDE},
{8'hE9, 8'hD0, 8'hD8},
{8'hD9, 8'hC0, 8'hC9},
{8'hE3, 8'hCE, 8'hD5},
{8'hF1, 8'hE3, 8'hE9},
{8'hFC, 8'hF5, 8'hF9},
{8'hFD, 8'hF9, 8'hFB},
{8'hF9, 8'hF6, 8'hF7},
{8'hED, 8'hEA, 8'hEC},
{8'hE2, 8'hD0, 8'hDA},
{8'hDD, 8'hC8, 8'hD2},
{8'hDD, 8'hC7, 8'hCE},
{8'hDE, 8'hC7, 8'hCE},
{8'hE6, 8'hD1, 8'hD8},
{8'hD6, 8'hC5, 8'hCE},
{8'hC0, 8'hB3, 8'hBF},
{8'hAD, 8'hA1, 8'hAF},
{8'h9C, 8'h83, 8'h97},
{8'h7E, 8'h71, 8'h93},
{8'h4F, 8'h5A, 8'h91},
{8'h29, 8'h4D, 8'h97},
{8'h1B, 8'h50, 8'hA5},
{8'h18, 8'h54, 8'hAF},
{8'h18, 8'h55, 8'hB0},
{8'h0F, 8'h40, 8'h97},
{8'h02, 8'h05, 8'h2B},
{8'h05, 8'h06, 8'h23},
{8'h00, 8'h02, 8'h18},
{8'h00, 8'h00, 8'h07},
{8'h6A, 8'h6A, 8'h65},
{8'hF3, 8'hEF, 8'hDA},
{8'hF4, 8'hE9, 8'hC5},
{8'hF3, 8'hE6, 8'hB8},
{8'hE0, 8'hE2, 8'hBC},
{8'hEF, 8'hF1, 8'hD1},
{8'hEE, 8'hED, 8'hD4},
{8'hE8, 8'hE6, 8'hD4},
{8'hFB, 8'hF9, 8'hEB},
{8'hF7, 8'hF4, 8'hE5},
{8'hE7, 8'hE0, 8'hCF},
{8'hFC, 8'hF6, 8'hE4},
{8'hE1, 8'hD6, 8'hCC},
{8'hF5, 8'hF0, 8'hE2},
{8'hFE, 8'hFC, 8'hE6},
{8'hED, 8'hE4, 8'hC8},
{8'hF7, 8'hE8, 8'hC6},
{8'hFD, 8'hF3, 8'hC7},
{8'hED, 8'hF5, 8'hBC},
{8'hE2, 8'hFB, 8'hBB},
{8'hF0, 8'hF0, 8'hC2},
{8'hF9, 8'hF4, 8'hCC},
{8'hE5, 8'hD9, 8'hB5},
{8'hDA, 8'hCC, 8'hAA},
{8'hC3, 8'hB5, 8'h92},
{8'hC7, 8'hBC, 8'h93},
{8'hF5, 8'hF1, 8'hC0},
{8'hF3, 8'hF3, 8'hBF},
{8'hDE, 8'hE0, 8'hC2},
{8'h80, 8'h81, 8'h74},
{8'h80, 8'h7D, 8'h83},
{8'h80, 8'h7D, 8'h88},
{8'h7F, 8'h7C, 8'h80},
{8'h7F, 8'h7E, 8'h7C},
{8'h7F, 8'h7D, 8'h7F},
{8'h7F, 8'h7C, 8'h84},
{8'h92, 8'h78, 8'h77},
{8'hD2, 8'hB7, 8'hB5},
{8'hE8, 8'hD0, 8'hCD},
{8'hDC, 8'hC1, 8'hBE},
{8'hC1, 8'hA5, 8'hA2},
{8'hB3, 8'h95, 8'h90},
{8'hAA, 8'h89, 8'h84},
{8'hA4, 8'h82, 8'h7C},
{8'hC5, 8'hA3, 8'h9C},
{8'hFC, 8'hE7, 8'hDE},
{8'hFF, 8'hED, 8'hE2},
{8'hFF, 8'hEC, 8'hDF},
{8'hF7, 8'hDE, 8'hCF},
{8'hE0, 8'hBE, 8'hAF},
{8'hEA, 8'hC6, 8'hB7},
{8'hFE, 8'hE5, 8'hD7},
{8'hF8, 8'hF4, 8'hEE},
{8'hFA, 8'hF6, 8'hF1},
{8'hFA, 8'hF1, 8'hEB},
{8'hFD, 8'hF2, 8'hE8},
{8'hFE, 8'hED, 8'hDC},
{8'hFB, 8'hDE, 8'hC6},
{8'hEF, 8'hC2, 8'hA4},
{8'hE6, 8'hAE, 8'h8A},
{8'hC0, 8'h82, 8'h67},
{8'h83, 8'h2C, 8'h3A},
{8'hE0, 8'h9F, 8'h6B},
{8'hB9, 8'hB7, 8'h7A},
{8'h23, 8'h56, 8'hAA},
{8'h0E, 8'h5A, 8'hBD},
{8'h18, 8'h3C, 8'h9C},
{8'h13, 8'h0B, 8'h45},
{8'h04, 8'h03, 8'h21},
{8'h00, 8'h00, 8'h1A},
{8'h00, 8'h00, 8'h0F},
{8'h1B, 8'h20, 8'h24},
{8'h5C, 8'h62, 8'h57},
{8'hA0, 8'hA7, 8'h8C},
{8'hBB, 8'hC3, 8'h9A},
{8'hCF, 8'hD6, 8'hA8},
{8'hEB, 8'hF2, 8'hC9},
{8'hF9, 8'hFF, 8'hD4},
{8'hEA, 8'hF5, 8'hC2},
{8'hEA, 8'hF3, 8'hC1},
{8'hE3, 8'hEB, 8'hC1},
{8'hE8, 8'hEE, 8'hD2},
{8'hF2, 8'hF6, 8'hE9},
{8'hF9, 8'hFB, 8'hF8},
{8'hED, 8'hF1, 8'hE2},
{8'hE4, 8'hE8, 8'hD2},
{8'hE6, 8'hE7, 8'hD0},
{8'hF0, 8'hF0, 8'hE1},
{8'hF6, 8'hF4, 8'hEF},
{8'hF2, 8'hEE, 8'hE7},
{8'hEC, 8'hE8, 8'hD3},
{8'hBA, 8'hB9, 8'h94},
{8'hD8, 8'hE1, 8'hA6},
{8'hE5, 8'hED, 8'hBC},
{8'hEA, 8'hED, 8'hD1},
{8'hF6, 8'hF7, 8'hEC},
{8'hFB, 8'hF9, 8'hF8},
{8'hF8, 8'hF4, 8'hF4},
{8'hF8, 8'hF5, 8'hF0},
{8'hFE, 8'hFB, 8'hF1},
{8'hF0, 8'hE9, 8'hDC},
{8'hFC, 8'hF6, 8'hE9},
{8'hF5, 8'hED, 8'hE2},
{8'hE9, 8'hE0, 8'hDA},
{8'hEE, 8'hE5, 8'hE5},
{8'hE6, 8'hDD, 8'hE4},
{8'h9A, 8'h90, 8'h9F},
{8'h96, 8'h8B, 8'h9C},
{8'hDD, 8'hCD, 8'hD3},
{8'hF7, 8'hEB, 8'hF0},
{8'hFF, 8'hF7, 8'hFC},
{8'hFF, 8'hFA, 8'hFE},
{8'hFD, 8'hFB, 8'hFD},
{8'hFC, 8'hFC, 8'hFD},
{8'hFD, 8'hFD, 8'hFD},
{8'hFE, 8'hFF, 8'hFF},
{8'hFE, 8'hF8, 8'hFD},
{8'hFA, 8'hEF, 8'hF5},
{8'hF0, 8'hE3, 8'hE9},
{8'hDB, 8'hCE, 8'hD7},
{8'h78, 8'h6F, 8'h7D},
{8'h1F, 8'h1D, 8'h32},
{8'h13, 8'h15, 8'h34},
{8'h06, 8'h0D, 8'h33},
{8'h00, 8'h0D, 8'h4E},
{8'h10, 8'h33, 8'h7B},
{8'h18, 8'h4F, 8'hA2},
{8'h0D, 8'h53, 8'hB4},
{8'h10, 8'h57, 8'hC0},
{8'h17, 8'h52, 8'hB4},
{8'h24, 8'h50, 8'hA0},
{8'h07, 8'h1C, 8'h5A},
{8'h01, 8'h01, 8'h20},
{8'h07, 8'h07, 8'h23},
{8'h00, 8'h01, 8'h14},
{8'h1E, 8'h1F, 8'h26},
{8'hD6, 8'hD6, 8'hC7},
{8'hEB, 8'hE8, 8'hCA},
{8'hE4, 8'hDC, 8'hB9},
{8'hE1, 8'hD6, 8'hB6},
{8'hEF, 8'hE6, 8'hD1},
{8'hF3, 8'hED, 8'hD9},
{8'hE4, 8'hDE, 8'hCB},
{8'hF5, 8'hEB, 8'hDB},
{8'hFF, 8'hF3, 8'hE8},
{8'hEF, 8'hE1, 8'hD8},
{8'hE5, 8'hD8, 8'hCD},
{8'hF0, 8'hEB, 8'hDF},
{8'hDB, 8'hD3, 8'hC8},
{8'hF7, 8'hF0, 8'hE2},
{8'hFF, 8'hFB, 8'hE7},
{8'hF2, 8'hEC, 8'hD0},
{8'hDE, 8'hD8, 8'hB4},
{8'hF4, 8'hF5, 8'hC7},
{8'hE7, 8'hF5, 8'hBD},
{8'hE2, 8'hF9, 8'hBB},
{8'hE7, 8'hF4, 8'hBF},
{8'hEB, 8'hF5, 8'hC2},
{8'hEE, 8'hF6, 8'hC5},
{8'hED, 8'hF3, 8'hC5},
{8'hEB, 8'hEE, 8'hC2},
{8'hEE, 8'hF3, 8'hC5},
{8'hEE, 8'hF5, 8'hC4},
{8'hF0, 8'hF8, 8'hC6},
{8'hEC, 8'hF0, 8'hCB},
{8'h9A, 8'h9B, 8'h8A},
{8'h78, 8'h76, 8'h79},
{8'h80, 8'h7C, 8'h88},
{8'h7F, 8'h7D, 8'h82},
{8'h7F, 8'h7D, 8'h7D},
{8'h7F, 8'h7D, 8'h7F},
{8'h7F, 8'h7D, 8'h82},
{8'h87, 8'h70, 8'h6E},
{8'h86, 8'h6F, 8'h6D},
{8'h8D, 8'h75, 8'h71},
{8'h8B, 8'h72, 8'h6E},
{8'h8A, 8'h70, 8'h6B},
{8'h85, 8'h6A, 8'h64},
{8'h99, 8'h7D, 8'h77},
{8'hBC, 8'hA2, 8'h9B},
{8'hE0, 8'hC9, 8'hBF},
{8'hEC, 8'hD8, 8'hCE},
{8'hED, 8'hD6, 8'hC9},
{8'hF2, 8'hE2, 8'hD4},
{8'hFE, 8'hEE, 8'hDF},
{8'hFF, 8'hEF, 8'hE0},
{8'hFF, 8'hEE, 8'hDF},
{8'hFF, 8'hE9, 8'hDD},
{8'hFB, 8'hF1, 8'hE9},
{8'hFD, 8'hF4, 8'hEC},
{8'hFF, 8'hF2, 8'hEB},
{8'hF7, 8'hE2, 8'hD7},
{8'hE1, 8'hC1, 8'hB2},
{8'hCB, 8'h9C, 8'h87},
{8'hA3, 8'h69, 8'h50},
{8'h78, 8'h3B, 8'h23},
{8'h3F, 8'h12, 8'h0D},
{8'h3C, 8'h09, 8'h11},
{8'hE6, 8'hC4, 8'h7E},
{8'h95, 8'h9D, 8'h73},
{8'h20, 8'h46, 8'hA6},
{8'h0F, 8'h40, 8'h99},
{8'h03, 8'h14, 8'h3F},
{8'h0B, 8'h00, 8'h1B},
{8'h01, 8'h03, 8'h14},
{8'h35, 8'h39, 8'h44},
{8'h89, 8'h91, 8'h91},
{8'hB2, 8'hBD, 8'hAE},
{8'hD5, 8'hE0, 8'hC1},
{8'hDA, 8'hE7, 8'hBB},
{8'hCF, 8'hDC, 8'hA6},
{8'hC4, 8'hD2, 8'h98},
{8'hDC, 8'hE4, 8'hCA},
{8'hF4, 8'hFB, 8'hE1},
{8'hEF, 8'hF6, 8'hD9},
{8'hE9, 8'hF0, 8'hD0},
{8'hE8, 8'hEE, 8'hCD},
{8'hE5, 8'hEC, 8'hCA},
{8'hE3, 8'hE9, 8'hC6},
{8'hE1, 8'hE7, 8'hC6},
{8'hED, 8'hE8, 8'hD9},
{8'hF0, 8'hEB, 8'hD9},
{8'hF5, 8'hF2, 8'hDE},
{8'hFC, 8'hF8, 8'hEC},
{8'hF9, 8'hF7, 8'hF2},
{8'hF6, 8'hF5, 8'hEB},
{8'hD4, 8'hD6, 8'hBB},
{8'hAA, 8'hB1, 8'h84},
{8'hB5, 8'hBF, 8'h89},
{8'hE7, 8'hF0, 8'hC4},
{8'hD9, 8'hDD, 8'hC3},
{8'hE9, 8'hE9, 8'hDF},
{8'hFE, 8'hFE, 8'hFB},
{8'hFD, 8'hFA, 8'hF6},
{8'hF8, 8'hF4, 8'hEB},
{8'hF9, 8'hF4, 8'hE5},
{8'hF7, 8'hF1, 8'hD0},
{8'hED, 8'hE6, 8'hC6},
{8'hEA, 8'hE5, 8'hC8},
{8'hE6, 8'hE0, 8'hCC},
{8'hEA, 8'hE4, 8'hDC},
{8'hF4, 8'hF0, 8'hF5},
{8'h2C, 8'h27, 8'h39},
{8'h0A, 8'h03, 8'h1C},
{8'h97, 8'h90, 8'h95},
{8'hBB, 8'hB6, 8'hB8},
{8'hBC, 8'hB7, 8'hB9},
{8'hB2, 8'hAF, 8'hB0},
{8'hA9, 8'hA7, 8'hA8},
{8'hA7, 8'hA6, 8'hA6},
{8'hA8, 8'hA9, 8'hA9},
{8'hAE, 8'hAF, 8'hAE},
{8'hB3, 8'hB2, 8'hB2},
{8'hB5, 8'hB3, 8'hB3},
{8'hD0, 8'hCF, 8'hD2},
{8'hBE, 8'hBD, 8'hCA},
{8'h19, 8'h1D, 8'h36},
{8'h08, 8'h11, 8'h3D},
{8'h0F, 8'h29, 8'h62},
{8'h17, 8'h3D, 8'h81},
{8'h19, 8'h4E, 8'hAD},
{8'h18, 8'h5A, 8'hB5},
{8'h05, 8'h53, 8'hAE},
{8'h06, 8'h58, 8'hBC},
{8'h10, 8'h56, 8'hC1},
{8'h24, 8'h53, 8'hB0},
{8'h18, 8'h2D, 8'h6D},
{8'h00, 8'h03, 8'h25},
{8'h01, 8'h02, 8'h17},
{8'h02, 8'h02, 8'h1D},
{8'h04, 8'h04, 8'h15},
{8'h9A, 8'h98, 8'h9C},
{8'hF8, 8'hF7, 8'hE0},
{8'hE0, 8'hDE, 8'hB8},
{8'hDD, 8'hD8, 8'hB8},
{8'hDB, 8'hD2, 8'hBE},
{8'hF8, 8'hE6, 8'hDD},
{8'hF6, 8'hEA, 8'hDD},
{8'hDF, 8'hD8, 8'hC5},
{8'hF8, 8'hE9, 8'hD8},
{8'hFF, 8'hED, 8'hE1},
{8'hEB, 8'hD4, 8'hCD},
{8'hC5, 8'hB5, 8'hAD},
{8'hEA, 8'hED, 8'hE2},
{8'hD8, 8'hD1, 8'hC2},
{8'hF4, 8'hE7, 8'hD8},
{8'hFF, 8'hF2, 8'hE0},
{8'hF7, 8'hED, 8'hD3},
{8'hDA, 8'hD8, 8'hB5},
{8'hEC, 8'hF4, 8'hC9},
{8'hE4, 8'hF1, 8'hC0},
{8'hE8, 8'hF6, 8'hC2},
{8'hE7, 8'hF9, 8'hC1},
{8'hE3, 8'hF6, 8'hBE},
{8'hE1, 8'hF4, 8'hBD},
{8'hE4, 8'hF4, 8'hC0},
{8'hE9, 8'hF7, 8'hC5},
{8'hE9, 8'hF5, 8'hC6},
{8'hE9, 8'hF3, 8'hC7},
{8'hEA, 8'hF3, 8'hC7},
{8'hF5, 8'hFA, 8'hD0},
{8'hB0, 8'hB2, 8'h9D},
{8'h7C, 8'h7A, 8'h7C},
{8'h7C, 8'h78, 8'h85},
{8'h7F, 8'h7C, 8'h84},
{8'h7F, 8'h7D, 8'h7F},
{8'h7F, 8'h7D, 8'h7E},
{8'h7F, 8'h7D, 8'h82},
{8'h89, 8'h82, 8'h7D},
{8'h85, 8'h7E, 8'h78},
{8'h82, 8'h7B, 8'h75},
{8'h83, 8'h7A, 8'h74},
{8'h89, 8'h80, 8'h77},
{8'hB6, 8'hAB, 8'hA2},
{8'hDC, 8'hD0, 8'hC6},
{8'hE1, 8'hD7, 8'hCC},
{8'hF5, 8'hE4, 8'hD9},
{8'hFC, 8'hEB, 8'hDF},
{8'hFB, 8'hEE, 8'hE0},
{8'hF1, 8'hE4, 8'hD6},
{8'hED, 8'hDA, 8'hCC},
{8'hFB, 8'hE9, 8'hDC},
{8'hF9, 8'hE6, 8'hDA},
{8'hFB, 8'hE4, 8'hD8},
{8'hFF, 8'hEB, 8'hD2},
{8'hFB, 8'hDD, 8'hC6},
{8'hE5, 8'hC3, 8'hAF},
{8'hC1, 8'h9C, 8'h8D},
{8'hA6, 8'h7E, 8'h73},
{8'h98, 8'h6D, 8'h63},
{8'h66, 8'h36, 8'h2D},
{8'h45, 8'h14, 8'h0C},
{8'h12, 8'h00, 8'h08},
{8'h3B, 8'h27, 8'h0D},
{8'hE4, 8'hDC, 8'h77},
{8'h7F, 8'h7C, 8'h70},
{8'h1A, 8'h27, 8'h59},
{8'h00, 8'h0A, 8'h47},
{8'h00, 8'h02, 8'h20},
{8'h02, 8'h05, 8'h01},
{8'h5F, 8'h66, 8'h58},
{8'hC1, 8'hC9, 8'hB8},
{8'hB3, 8'hBA, 8'hA5},
{8'hB1, 8'hB7, 8'h9C},
{8'hBB, 8'hC2, 8'hA2},
{8'hBE, 8'hC6, 8'hA3},
{8'hAD, 8'hB9, 8'h93},
{8'hDC, 8'hE8, 8'hC2},
{8'hE7, 8'hEC, 8'hD1},
{8'hF2, 8'hF4, 8'hDE},
{8'hFD, 8'hFE, 8'hEC},
{8'hF6, 8'hF7, 8'hE7},
{8'hF4, 8'hF3, 8'hDF},
{8'hF0, 8'hF0, 8'hD3},
{8'hEA, 8'hEA, 8'hC4},
{8'hE6, 8'hE7, 8'hB9},
{8'hF2, 8'hEA, 8'hC4},
{8'hFC, 8'hF5, 8'hD1},
{8'hFE, 8'hFB, 8'hDC},
{8'hFE, 8'hFB, 8'hE6},
{8'hF4, 8'hF2, 8'hE9},
{8'hDF, 8'hE1, 8'hD6},
{8'hBA, 8'hC3, 8'hA7},
{8'hAA, 8'hB6, 8'h89},
{8'hB4, 8'hBF, 8'h8F},
{8'hD1, 8'hD9, 8'hB4},
{8'h8D, 8'h91, 8'h7C},
{8'h9D, 8'h9D, 8'h95},
{8'hDE, 8'hDB, 8'hD8},
{8'hFD, 8'hFC, 8'hF3},
{8'hF3, 8'hEE, 8'hDE},
{8'hEA, 8'hE5, 8'hCC},
{8'hEA, 8'hE6, 8'hA7},
{8'hD5, 8'hD1, 8'h93},
{8'hE1, 8'hDF, 8'hA7},
{8'hE7, 8'hE5, 8'hB9},
{8'hE5, 8'hE4, 8'hCA},
{8'hC7, 8'hC6, 8'hC1},
{8'h3C, 8'h39, 8'h47},
{8'h2A, 8'h28, 8'h3E},
{8'hB1, 8'hB2, 8'hB4},
{8'hD1, 8'hD2, 8'hD2},
{8'hE2, 8'hE3, 8'hE2},
{8'hEF, 8'hEF, 8'hEF},
{8'hF5, 8'hF5, 8'hF5},
{8'hF8, 8'hF7, 8'hF8},
{8'hF5, 8'hF4, 8'hF5},
{8'hEE, 8'hED, 8'hED},
{8'hDE, 8'hE1, 8'hDC},
{8'hCA, 8'hCE, 8'hCC},
{8'hBD, 8'hC0, 8'hC2},
{8'h5F, 8'h66, 8'h76},
{8'h1D, 8'h31, 8'h56},
{8'h39, 8'h5E, 8'h9C},
{8'h21, 8'h55, 8'hA6},
{8'h1A, 8'h57, 8'hB4},
{8'h14, 8'h51, 8'hB6},
{8'h0F, 8'h54, 8'hAC},
{8'h0F, 8'h5C, 8'hAA},
{8'h0D, 8'h58, 8'hAE},
{8'h14, 8'h4F, 8'hB0},
{8'h1E, 8'h3E, 8'h94},
{8'h02, 8'h07, 8'h38},
{8'h06, 8'h02, 8'h12},
{8'h01, 8'h03, 8'h13},
{8'h00, 8'h00, 8'h18},
{8'h3E, 8'h3D, 8'h57},
{8'hEF, 8'hED, 8'hEE},
{8'hDE, 8'hDD, 8'hBF},
{8'hC1, 8'hC0, 8'h94},
{8'hD8, 8'hD5, 8'hB6},
{8'hEC, 8'hE4, 8'hD9},
{8'hF3, 8'hE1, 8'hDC},
{8'hF8, 8'hF0, 8'hE3},
{8'hE0, 8'hDD, 8'hC8},
{8'hF1, 8'hE0, 8'hCB},
{8'hFF, 8'hE9, 8'hDB},
{8'hF3, 8'hDA, 8'hD1},
{8'hBB, 8'hAF, 8'hA6},
{8'hDC, 8'hE8, 8'hDC},
{8'hE5, 8'hDB, 8'hC8},
{8'hEA, 8'hD8, 8'hC6},
{8'hFF, 8'hEE, 8'hDC},
{8'hFB, 8'hED, 8'hD3},
{8'hD3, 8'hD3, 8'hB2},
{8'hDF, 8'hEA, 8'hC1},
{8'hE5, 8'hEF, 8'hC4},
{8'hEF, 8'hF4, 8'hC9},
{8'hE5, 8'hF4, 8'hBE},
{8'hEA, 8'hFB, 8'hC4},
{8'hED, 8'hFE, 8'hC7},
{8'hEA, 8'hF9, 8'hC3},
{8'hEB, 8'hF8, 8'hC6},
{8'hED, 8'hF5, 8'hCA},
{8'hED, 8'hF0, 8'hCB},
{8'hEA, 8'hEB, 8'hC8},
{8'hF1, 8'hF7, 8'hC8},
{8'hA8, 8'hAA, 8'h90},
{8'h79, 8'h77, 8'h79},
{8'h80, 8'h7C, 8'h8A},
{8'h80, 8'h7C, 8'h86},
{8'h7F, 8'h7D, 8'h7F},
{8'h7F, 8'h7D, 8'h7E},
{8'h7F, 8'h7D, 8'h81},
{8'h7C, 8'h81, 8'h7E},
{8'h7B, 8'h7F, 8'h7A},
{8'h7C, 8'h7A, 8'h72},
{8'hA8, 8'hA5, 8'h99},
{8'hE6, 8'hE2, 8'hD5},
{8'hF6, 8'hF0, 8'hE3},
{8'hE9, 8'hE4, 8'hD9},
{8'hD4, 8'hD0, 8'hC4},
{8'hE2, 8'hCC, 8'hBD},
{8'hD3, 8'hBA, 8'hA9},
{8'hD4, 8'hB6, 8'hA6},
{8'hEA, 8'hCD, 8'hBC},
{8'hFD, 8'hE7, 8'hD6},
{8'hFF, 8'hE8, 8'hD8},
{8'hF9, 8'hDB, 8'hCC},
{8'hE2, 8'hBF, 8'hAF},
{8'hCF, 8'hA6, 8'h8D},
{8'hB4, 8'h8B, 8'h75},
{8'h95, 8'h73, 8'h64},
{8'h8F, 8'h74, 8'h6D},
{8'h91, 8'h78, 8'h76},
{8'h95, 8'h79, 8'h79},
{8'h74, 8'h54, 8'h53},
{8'h3C, 8'h19, 8'h1A},
{8'h1C, 8'h04, 8'h1B},
{8'h5D, 8'h51, 8'h1E},
{8'hDE, 8'hD9, 8'h7A},
{8'h43, 8'h38, 8'h43},
{8'h05, 8'h05, 8'h15},
{8'h00, 8'h01, 8'h15},
{8'h0B, 8'h0E, 8'h1B},
{8'h5C, 8'h69, 8'h50},
{8'h92, 8'h99, 8'h85},
{8'h7E, 8'h84, 8'h70},
{8'h6F, 8'h73, 8'h5E},
{8'hA4, 8'hA8, 8'h90},
{8'hC5, 8'hCA, 8'hAF},
{8'hA7, 8'hAF, 8'h8F},
{8'hBF, 8'hC8, 8'hA7},
{8'hEB, 8'hF6, 8'hD2},
{8'hE5, 8'hEE, 8'hC1},
{8'hEA, 8'hF1, 8'hCC},
{8'hF7, 8'hF8, 8'hE2},
{8'hFB, 8'hF9, 8'hED},
{8'hF4, 8'hEF, 8'hE2},
{8'hF5, 8'hEF, 8'hD8},
{8'hF4, 8'hEF, 8'hCA},
{8'hF2, 8'hED, 8'hBE},
{8'hF8, 8'hEA, 8'hAB},
{8'hEB, 8'hDE, 8'h8B},
{8'hEA, 8'hE3, 8'h90},
{8'hF9, 8'hF3, 8'hC1},
{8'hF9, 8'hF3, 8'hE0},
{8'hC8, 8'hC8, 8'hB8},
{8'hBA, 8'hC0, 8'hA6},
{8'hBF, 8'hC9, 8'hAA},
{8'hB3, 8'hBA, 8'hA1},
{8'hD1, 8'hD5, 8'hC1},
{8'hC8, 8'hC8, 8'hBC},
{8'hD7, 8'hD5, 8'hD1},
{8'hF0, 8'hEB, 8'hEB},
{8'hF7, 8'hF2, 8'hEC},
{8'hF3, 8'hEE, 8'hDC},
{8'hEE, 8'hEA, 8'hC9},
{8'hDA, 8'hD7, 8'h87},
{8'hBB, 8'hB8, 8'h68},
{8'hD4, 8'hD3, 8'h8B},
{8'hE2, 8'hE1, 8'hA9},
{8'hF1, 8'hF1, 8'hCD},
{8'h98, 8'h98, 8'h8B},
{8'h57, 8'h56, 8'h5F},
{8'h6E, 8'h6E, 8'h80},
{8'hFE, 8'hFF, 8'hFF},
{8'hFF, 8'hFF, 8'hFF},
{8'hFB, 8'hFC, 8'hFC},
{8'hFB, 8'hFC, 8'hFC},
{8'hFD, 8'hFD, 8'hFD},
{8'hFE, 8'hFD, 8'hFE},
{8'hFF, 8'hFF, 8'hFF},
{8'hFF, 8'hFF, 8'hFF},
{8'hFC, 8'hFF, 8'hFF},
{8'hFF, 8'hFF, 8'hFF},
{8'hF3, 8'hF5, 8'hFA},
{8'h53, 8'h62, 8'h7F},
{8'h4C, 8'h5E, 8'h86},
{8'h67, 8'h84, 8'hBF},
{8'h1F, 8'h55, 8'hAF},
{8'h12, 8'h53, 8'hBD},
{8'h19, 8'h4F, 8'hB1},
{8'h13, 8'h53, 8'hAC},
{8'h13, 8'h5B, 8'hAF},
{8'h19, 8'h5A, 8'hAC},
{8'h22, 8'h4C, 8'h9B},
{8'h09, 8'h13, 8'h52},
{8'h04, 8'h00, 8'h21},
{8'h0C, 8'h04, 8'h15},
{8'h03, 8'h02, 8'h18},
{8'h0A, 8'h08, 8'h1E},
{8'hBA, 8'hB7, 8'hBF},
{8'hDF, 8'hDD, 8'hD2},
{8'hAD, 8'hAB, 8'h8E},
{8'hBF, 8'hBC, 8'h9C},
{8'hD6, 8'hD1, 8'hC0},
{8'hEB, 8'hE4, 8'hE2},
{8'hF3, 8'hE7, 8'hE8},
{8'hF8, 8'hF2, 8'hEA},
{8'hE9, 8'hE5, 8'hD1},
{8'hE5, 8'hD3, 8'hBC},
{8'hFD, 8'hE3, 8'hD2},
{8'hE8, 8'hCE, 8'hC1},
{8'hC7, 8'hBD, 8'hAD},
{8'hCD, 8'hD7, 8'hC2},
{8'hF1, 8'hE6, 8'hDA},
{8'hDA, 8'hCB, 8'hBD},
{8'hFA, 8'hE5, 8'hD3},
{8'hFD, 8'hE8, 8'hD1},
{8'hD0, 8'hC3, 8'hA9},
{8'hE3, 8'hE2, 8'hC4},
{8'hF0, 8'hF3, 8'hD0},
{8'hEC, 8'hEF, 8'hC8},
{8'hEA, 8'hF4, 8'hBD},
{8'hEE, 8'hF8, 8'hC4},
{8'hCB, 8'hD5, 8'hA6},
{8'hAA, 8'hB1, 8'h8E},
{8'hA2, 8'hA7, 8'h8D},
{8'h98, 8'h9A, 8'h85},
{8'h91, 8'h90, 8'h77},
{8'hAC, 8'hAB, 8'h8D},
{8'hD5, 8'hD8, 8'hB9},
{8'h84, 8'h86, 8'h75},
{8'h80, 8'h7E, 8'h7F},
{8'h81, 8'h7E, 8'h87},
{8'h7E, 8'h7B, 8'h82},
{8'h7F, 8'h7D, 8'h7F},
{8'h7F, 8'h7D, 8'h7E},
{8'h7F, 8'h7D, 8'h7F},
{8'h82, 8'h78, 8'h7D},
{8'h8C, 8'h7C, 8'h7C},
{8'hD7, 8'hBD, 8'hB5},
{8'hFF, 8'hEE, 8'hDF},
{8'hFA, 8'hDE, 8'hCD},
{8'hF3, 8'hDA, 8'hCC},
{8'hF9, 8'hE4, 8'hDC},
{8'hF4, 8'hE2, 8'hDD},
{8'hE6, 8'hC2, 8'hB2},
{8'hCA, 8'hA0, 8'h90},
{8'hA4, 8'h76, 8'h66},
{8'h97, 8'h69, 8'h59},
{8'hAE, 8'h85, 8'h75},
{8'hC7, 8'h9D, 8'h8D},
{8'hC3, 8'h98, 8'h88},
{8'hA5, 8'h7A, 8'h6B},
{8'h89, 8'h72, 8'h6B},
{8'h87, 8'h77, 8'h76},
{8'h81, 8'h7A, 8'h80},
{8'h7B, 8'h7B, 8'h85},
{8'h7E, 8'h7E, 8'h88},
{8'h82, 8'h7B, 8'h81},
{8'h7C, 8'h6D, 8'h6A},
{8'h41, 8'h27, 8'h22},
{8'h4A, 8'h08, 8'h0B},
{8'h89, 8'h5B, 8'h30},
{8'h90, 8'h77, 8'h43},
{8'h09, 8'h00, 8'h0B},
{8'h00, 8'h00, 8'h10},
{8'h24, 8'h2F, 8'h18},
{8'hAA, 8'hB5, 8'h84},
{8'hE1, 8'hE4, 8'hD1},
{8'h8D, 8'h92, 8'h8F},
{8'h81, 8'h86, 8'h81},
{8'h7C, 8'h82, 8'h7A},
{8'hB9, 8'hC0, 8'hB0},
{8'hC0, 8'hC9, 8'hAE},
{8'hA3, 8'hAE, 8'h87},
{8'hE3, 8'hF0, 8'hBC},
{8'hE7, 8'hF5, 8'hBA},
{8'hE2, 8'hF2, 8'hB9},
{8'hE4, 8'hF1, 8'hC4},
{8'hEE, 8'hF4, 8'hDA},
{8'hFC, 8'hFC, 8'hEE},
{8'hFA, 8'hF7, 8'hE9},
{8'hF7, 8'hF4, 8'hDA},
{8'hF6, 8'hF3, 8'hC9},
{8'hF8, 8'hF4, 8'hC0},
{8'hF8, 8'hE1, 8'h99},
{8'hEA, 8'hD9, 8'h58},
{8'hDE, 8'hD5, 8'h44},
{8'hE0, 8'hD5, 8'h80},
{8'hEF, 8'hE2, 8'hC3},
{8'hEA, 8'hE4, 8'hCC},
{8'hC3, 8'hC2, 8'hA8},
{8'hE3, 8'hE3, 8'hD9},
{8'hEC, 8'hE9, 8'hEF},
{8'hF5, 8'hF2, 8'hF2},
{8'hFC, 8'hF8, 8'hF2},
{8'hF9, 8'hF4, 8'hF2},
{8'hF9, 8'hF2, 8'hF7},
{8'hFA, 8'hF1, 8'hF2},
{8'hEF, 8'hEA, 8'hD9},
{8'hE7, 8'hE2, 8'hBF},
{8'hDD, 8'hD6, 8'h90},
{8'hCC, 8'hC7, 8'h80},
{8'hE5, 8'hE2, 8'hA4},
{8'hDD, 8'hDA, 8'hAA},
{8'hEE, 8'hEB, 8'hCE},
{8'h6F, 8'h6D, 8'h67},
{8'h26, 8'h25, 8'h30},
{8'h55, 8'h52, 8'h69},
{8'hC7, 8'hC3, 8'hC6},
{8'hDB, 8'hD3, 8'hD6},
{8'hF7, 8'hF2, 8'hF4},
{8'hFF, 8'hFF, 8'hFF},
{8'hFF, 8'hFF, 8'hFF},
{8'hF6, 8'hF6, 8'hF6},
{8'hE8, 8'hEB, 8'hE9},
{8'hDA, 8'hE1, 8'hE1},
{8'hC2, 8'hD5, 8'hD8},
{8'hCC, 8'hC1, 8'hB3},
{8'h8F, 8'h87, 8'h9D},
{8'h18, 8'h33, 8'h72},
{8'h45, 8'h56, 8'h87},
{8'h54, 8'h63, 8'h96},
{8'h1F, 8'h4F, 8'hA8},
{8'h19, 8'h51, 8'hBC},
{8'h1D, 8'h51, 8'hAF},
{8'h10, 8'h52, 8'hB9},
{8'h0B, 8'h55, 8'hBF},
{8'h1A, 8'h51, 8'hA9},
{8'h0C, 8'h1C, 8'h53},
{8'h05, 8'h00, 8'h1D},
{8'h09, 8'h00, 8'h15},
{8'h05, 8'h00, 8'h1B},
{8'h02, 8'h00, 8'h19},
{8'h71, 8'h6A, 8'h72},
{8'hE5, 8'hE2, 8'hCB},
{8'hD0, 8'hD0, 8'hAC},
{8'hA1, 8'hA0, 8'h85},
{8'hBC, 8'hB7, 8'hAD},
{8'hBC, 8'hB6, 8'hB4},
{8'hE7, 8'hE2, 8'hE3},
{8'hF3, 8'hF3, 8'hFB},
{8'hFB, 8'hF6, 8'hF4},
{8'hFD, 8'hF7, 8'hE4},
{8'hDF, 8'hC9, 8'hB3},
{8'hD7, 8'hBE, 8'hAE},
{8'hD5, 8'hC0, 8'hB1},
{8'hE3, 8'hD6, 8'hBC},
{8'hE4, 8'hDE, 8'hBD},
{8'hFD, 8'hF7, 8'hFB},
{8'hE6, 8'hDA, 8'hD6},
{8'hE5, 8'hCD, 8'hBD},
{8'hFB, 8'hDC, 8'hCC},
{8'hCD, 8'hAE, 8'hA3},
{8'hF2, 8'hE6, 8'hDA},
{8'hF0, 8'hEC, 8'hD3},
{8'hEB, 8'hF2, 8'hCA},
{8'hEA, 8'hF4, 8'hB9},
{8'hEF, 8'hF7, 8'hC2},
{8'hCC, 8'hD2, 8'hAE},
{8'h80, 8'h81, 8'h79},
{8'h76, 8'h74, 8'h81},
{8'h78, 8'h76, 8'h83},
{8'h77, 8'h79, 8'h71},
{8'h85, 8'h89, 8'h70},
{8'h82, 8'h80, 8'h81},
{8'h7B, 8'h79, 8'h7B},
{8'h7E, 8'h7C, 8'h7C},
{8'h7F, 8'h7D, 8'h7D},
{8'h7F, 8'h7D, 8'h7E},
{8'h7F, 8'h7D, 8'h7E},
{8'h7F, 8'h7D, 8'h7E},
{8'h7F, 8'h7D, 8'h7E},
{8'h94, 8'h6C, 8'h6D},
{8'hB2, 8'h84, 8'h81},
{8'hEC, 8'hB8, 8'hAE},
{8'hE4, 8'hAE, 8'hA0},
{8'hF5, 8'hC8, 8'hBA},
{8'hF5, 8'hC9, 8'hC0},
{8'hD1, 8'hA4, 8'hA0},
{8'hA5, 8'h7D, 8'h7C},
{8'h89, 8'h72, 8'h6E},
{8'h87, 8'h72, 8'h6D},
{8'h87, 8'h72, 8'h6D},
{8'h8E, 8'h79, 8'h75},
{8'h85, 8'h70, 8'h6B},
{8'h84, 8'h6E, 8'h6A},
{8'h85, 8'h70, 8'h6C},
{8'h87, 8'h72, 8'h6E},
{8'h88, 8'h77, 8'h70},
{8'h8C, 8'h80, 8'h7E},
{8'h7C, 8'h78, 8'h7B},
{8'h7D, 8'h7D, 8'h84},
{8'h7B, 8'h7C, 8'h83},
{8'h82, 8'h7E, 8'h81},
{8'h86, 8'h7B, 8'h78},
{8'h50, 8'h3A, 8'h35},
{8'h60, 8'h0C, 8'h0A},
{8'h98, 8'h55, 8'h1F},
{8'h65, 8'h3E, 8'h0F},
{8'h14, 8'h06, 8'h09},
{8'h69, 8'h67, 8'h6E},
{8'hD5, 8'hE0, 8'hB8},
{8'hEA, 8'hFB, 8'hBF},
{8'hE4, 8'hF3, 8'hD2},
{8'hB6, 8'hBD, 8'hA9},
{8'h89, 8'h90, 8'h7B},
{8'h88, 8'h90, 8'h7A},
{8'hD4, 8'hDD, 8'hC3},
{8'hB1, 8'hBB, 8'h9A},
{8'hC1, 8'hCC, 8'hA2},
{8'hEA, 8'hF6, 8'hC3},
{8'hE0, 8'hEE, 8'hB4},
{8'hE0, 8'hF0, 8'hB7},
{8'hE7, 8'hF2, 8'hC6},
{8'hD4, 8'hDA, 8'hBD},
{8'hE3, 8'hE5, 8'hD5},
{8'hEE, 8'hEC, 8'hDF},
{8'hF4, 8'hF1, 8'hDC},
{8'hF7, 8'hF3, 8'hD3},
{8'hF9, 8'hF3, 8'hCD},
{8'hFA, 8'hE8, 8'hB5},
{8'hEB, 8'hE0, 8'h7D},
{8'hDC, 8'hD7, 8'h68},
{8'hD9, 8'hD2, 8'h8F},
{8'hE7, 8'hDE, 8'hC4},
{8'hF2, 8'hEC, 8'hD7},
{8'hE7, 8'hE6, 8'hCD},
{8'hEE, 8'hEE, 8'hDC},
{8'hF6, 8'hF6, 8'hEC},
{8'hF3, 8'hF5, 8'hE3},
{8'hF9, 8'hF9, 8'hE4},
{8'hF9, 8'hF7, 8'hE8},
{8'hF7, 8'hF2, 8'hEE},
{8'hF7, 8'hF1, 8'hED},
{8'hEC, 8'hE7, 8'hD5},
{8'hE3, 8'hDF, 8'hBF},
{8'hE2, 8'hDB, 8'hAA},
{8'hDB, 8'hD4, 8'hA6},
{8'hEE, 8'hE8, 8'hC1},
{8'hEA, 8'hE6, 8'hCA},
{8'hCC, 8'hC8, 8'hBD},
{8'h32, 8'h2F, 8'h35},
{8'h00, 8'h00, 8'h0B},
{8'h7C, 8'h76, 8'h8F},
{8'hC5, 8'hBD, 8'hC0},
{8'h91, 8'h8B, 8'h8D},
{8'h73, 8'h6E, 8'h70},
{8'h8F, 8'h8B, 8'h8C},
{8'h75, 8'h73, 8'h74},
{8'h6E, 8'h6F, 8'h6E},
{8'h95, 8'h97, 8'h96},
{8'hB7, 8'hBB, 8'hBB},
{8'hBE, 8'hC1, 8'hC5},
{8'hB7, 8'h9F, 8'hA0},
{8'h4D, 8'h57, 8'h84},
{8'h0C, 8'h45, 8'h9F},
{8'h11, 8'h48, 8'h98},
{8'h1F, 8'h4F, 8'h9B},
{8'h17, 8'h53, 8'hB2},
{8'h17, 8'h51, 8'hB7},
{8'h1B, 8'h55, 8'hB6},
{8'h14, 8'h55, 8'hB8},
{8'h15, 8'h53, 8'hB2},
{8'h0A, 8'h2F, 8'h78},
{8'h00, 8'h01, 8'h30},
{8'h05, 8'h00, 8'h1A},
{8'h06, 8'h02, 8'h19},
{8'h04, 8'h03, 8'h1D},
{8'h26, 8'h21, 8'h28},
{8'hD5, 8'hD1, 8'hC4},
{8'hBB, 8'hBA, 8'h99},
{8'h93, 8'h93, 8'h6D},
{8'h99, 8'h98, 8'h7A},
{8'hA5, 8'hA3, 8'h8E},
{8'hD4, 8'hD1, 8'hBD},
{8'hE9, 8'hE8, 8'hD3},
{8'hF4, 8'hF4, 8'hF2},
{8'hFA, 8'hF7, 8'hEB},
{8'hF4, 8'hEB, 8'hD2},
{8'hE7, 8'hD5, 8'hBD},
{8'hC5, 8'hAE, 8'h9E},
{8'hF3, 8'hE2, 8'hD4},
{8'hE6, 8'hDB, 8'hC4},
{8'hE7, 8'hE3, 8'hC5},
{8'hFD, 8'hFB, 8'hF7},
{8'hFC, 8'hF6, 8'hEF},
{8'hD2, 8'hC0, 8'hB4},
{8'hB7, 8'h9B, 8'h94},
{8'hC0, 8'hA7, 8'hA5},
{8'hEF, 8'hE2, 8'hDA},
{8'hE6, 8'hE6, 8'hCB},
{8'hE5, 8'hF0, 8'hC4},
{8'hEA, 8'hF4, 8'hC0},
{8'hF1, 8'hF8, 8'hC5},
{8'hF1, 8'hF6, 8'hCA},
{8'hC3, 8'hC7, 8'hAE},
{8'hA2, 8'hA2, 8'h9E},
{8'h96, 8'h95, 8'h9A},
{8'h95, 8'h96, 8'h94},
{8'h89, 8'h8B, 8'h7F},
{8'h83, 8'h82, 8'h81},
{8'h89, 8'h87, 8'h89},
{8'h7E, 8'h7C, 8'h7D},
{8'h7D, 8'h7B, 8'h7C},
{8'h7F, 8'h7D, 8'h7E},
{8'h7F, 8'h7D, 8'h7E},
{8'h7F, 8'h7D, 8'h7E},
{8'h7F, 8'h7D, 8'h7E},
{8'h8E, 8'h6C, 8'h64},
{8'h93, 8'h6E, 8'h63},
{8'h8D, 8'h64, 8'h56},
{8'hA6, 8'h7B, 8'h6B},
{8'hAE, 8'h84, 8'h74},
{8'h95, 8'h70, 8'h66},
{8'h8F, 8'h71, 8'h6C},
{8'h8F, 8'h78, 8'h76},
{8'h82, 8'h7D, 8'h82},
{8'h80, 8'h7D, 8'h82},
{8'h80, 8'h7D, 8'h83},
{8'h81, 8'h7E, 8'h83},
{8'h80, 8'h7D, 8'h82},
{8'h82, 8'h7F, 8'h84},
{8'h80, 8'h7D, 8'h83},
{8'h7B, 8'h78, 8'h7D},
{8'h85, 8'h7B, 8'h76},
{8'h83, 8'h7D, 8'h7A},
{8'h83, 8'h82, 8'h85},
{8'h79, 8'h7C, 8'h81},
{8'h7A, 8'h7D, 8'h83},
{8'h7D, 8'h7D, 8'h7F},
{8'h85, 8'h80, 8'h7E},
{8'h68, 8'h58, 8'h54},
{8'h67, 8'h19, 8'h0F},
{8'h96, 8'h57, 8'h20},
{8'h79, 8'h55, 8'h27},
{8'hB8, 8'hA5, 8'h99},
{8'hEE, 8'hED, 8'hE2},
{8'hE6, 8'hF7, 8'hC2},
{8'hE0, 8'hF6, 8'hB1},
{8'hDF, 8'hF2, 8'hC3},
{8'hDA, 8'hE5, 8'hBC},
{8'hBE, 8'hC9, 8'hA1},
{8'hA3, 8'hAE, 8'h88},
{8'hDB, 8'hE5, 8'hBF},
{8'hB7, 8'hC2, 8'h99},
{8'hBD, 8'hC9, 8'h9A},
{8'hDF, 8'hEC, 8'hB6},
{8'hE8, 8'hF5, 8'hBC},
{8'hE2, 8'hEF, 8'hB8},
{8'hA6, 8'hB0, 8'h83},
{8'h8F, 8'h95, 8'h75},
{8'hD6, 8'hD8, 8'hC5},
{8'hE9, 8'hE7, 8'hDB},
{8'hFA, 8'hF6, 8'hE8},
{8'hFE, 8'hF9, 8'hE6},
{8'hF4, 8'hEE, 8'hD7},
{8'hF5, 8'hEC, 8'hCE},
{8'hEE, 8'hEA, 8'hAD},
{8'hE8, 8'hE7, 8'h9E},
{8'hE8, 8'hE5, 8'hB5},
{8'hF8, 8'hF3, 8'hDE},
{8'hEF, 8'hEC, 8'hDA},
{8'hEA, 8'hE8, 8'hCF},
{8'hEB, 8'hEA, 8'hD0},
{8'hE1, 8'hE4, 8'hC8},
{8'hD6, 8'hDB, 8'hB7},
{8'hCC, 8'hD0, 8'hA9},
{8'hE0, 8'hE1, 8'hC4},
{8'hF0, 8'hED, 8'hDE},
{8'hED, 8'hE9, 8'hDE},
{8'hEF, 8'hEB, 8'hD9},
{8'hE4, 8'hE0, 8'hC3},
{8'hDE, 8'hD6, 8'hB8},
{8'hE2, 8'hDB, 8'hC0},
{8'hED, 8'hE6, 8'hD2},
{8'hEC, 8'hE6, 8'hDB},
{8'hD5, 8'hCF, 8'hD0},
{8'h25, 8'h20, 8'h2E},
{8'h0A, 8'h06, 8'h1F},
{8'h79, 8'h74, 8'h8D},
{8'hA2, 8'h9D, 8'h9F},
{8'h9C, 8'h97, 8'h98},
{8'hB0, 8'hAD, 8'hAE},
{8'hC9, 8'hC7, 8'hC8},
{8'hC2, 8'hC1, 8'hC2},
{8'hA2, 8'hA1, 8'hA1},
{8'hA3, 8'hA3, 8'hA3},
{8'hB6, 8'hB5, 8'hB6},
{8'hCA, 8'hC0, 8'hC5},
{8'hCE, 8'hBE, 8'hD2},
{8'h42, 8'h59, 8'h9A},
{8'h10, 8'h53, 8'hBA},
{8'h0C, 8'h58, 8'hBB},
{8'h0F, 8'h57, 8'hB3},
{8'h0E, 8'h56, 8'hB9},
{8'h10, 8'h52, 8'hB9},
{8'h13, 8'h53, 8'hB6},
{8'h18, 8'h53, 8'hB0},
{8'h17, 8'h43, 8'h92},
{8'h01, 8'h0B, 8'h41},
{8'h03, 8'h01, 8'h20},
{8'h09, 8'h02, 8'h18},
{8'h04, 8'h02, 8'h1A},
{8'h01, 8'h03, 8'h18},
{8'h9A, 8'h99, 8'h88},
{8'hDB, 8'hD9, 8'hBC},
{8'h96, 8'h96, 8'h71},
{8'hAF, 8'hAF, 8'h8F},
{8'h92, 8'h90, 8'h79},
{8'hA0, 8'h9D, 8'h89},
{8'hDA, 8'hD9, 8'hBB},
{8'hE1, 8'hE2, 8'hBC},
{8'hEC, 8'hEB, 8'hDE},
{8'hFC, 8'hF9, 8'hE5},
{8'hE8, 8'hDF, 8'hC1},
{8'hDD, 8'hCC, 8'hB2},
{8'hEE, 8'hDB, 8'hCC},
{8'hFD, 8'hF0, 8'hE4},
{8'hEF, 8'hE6, 8'hD4},
{8'hE2, 8'hDF, 8'hC4},
{8'hF8, 8'hFA, 8'hEE},
{8'hF3, 8'hF2, 8'hE6},
{8'hFC, 8'hF4, 8'hEA},
{8'hE5, 8'hD3, 8'hD3},
{8'hE6, 8'hD2, 8'hD9},
{8'hE7, 8'hDE, 8'hD9},
{8'hED, 8'hF1, 8'hD5},
{8'hDC, 8'hEB, 8'hBB},
{8'hE9, 8'hF1, 8'hC8},
{8'hE9, 8'hF2, 8'hC1},
{8'hED, 8'hF6, 8'hBF},
{8'hD1, 8'hD9, 8'hAD},
{8'h88, 8'h8B, 8'h76},
{8'h89, 8'h89, 8'h87},
{8'h8F, 8'h8E, 8'h94},
{8'h92, 8'h92, 8'h95},
{8'h8D, 8'h8C, 8'h8D},
{8'h85, 8'h83, 8'h84},
{8'h7F, 8'h7D, 8'h7E},
{8'h80, 8'h7E, 8'h7F},
{8'h7F, 8'h7D, 8'h7E},
{8'h7F, 8'h7D, 8'h7E},
{8'h7F, 8'h7D, 8'h7E},
{8'h7F, 8'h7D, 8'h7E},
{8'h83, 8'h7D, 8'h72},
{8'h7B, 8'h73, 8'h67},
{8'h85, 8'h7B, 8'h6E},
{8'h7D, 8'h74, 8'h67},
{8'h80, 8'h7A, 8'h6F},
{8'h80, 8'h7F, 8'h77},
{8'h79, 8'h7D, 8'h7A},
{8'h77, 8'h7E, 8'h7F},
{8'h7B, 8'h7D, 8'h82},
{8'h7D, 8'h7F, 8'h84},
{8'h7C, 8'h7D, 8'h83},
{8'h7B, 8'h7D, 8'h82},
{8'h7C, 8'h7E, 8'h83},
{8'h7D, 8'h7E, 8'h84},
{8'h7D, 8'h7F, 8'h84},
{8'h7D, 8'h7E, 8'h83},
{8'h82, 8'h7E, 8'h7A},
{8'h81, 8'h7E, 8'h7C},
{8'h7F, 8'h80, 8'h81},
{8'h7B, 8'h7F, 8'h83},
{8'h7B, 8'h80, 8'h83},
{8'h7D, 8'h7E, 8'h7F},
{8'h81, 8'h7F, 8'h7E},
{8'h74, 8'h6C, 8'h68},
{8'h5E, 8'h38, 8'h21},
{8'hB3, 8'h99, 8'h5D},
{8'hEE, 8'hE5, 8'hA0},
{8'hF1, 8'hF2, 8'hCA},
{8'hE5, 8'hF0, 8'hCF},
{8'hDF, 8'hF1, 8'hB7},
{8'hE5, 8'hF9, 8'hB2},
{8'hE3, 8'hF2, 8'hB8},
{8'hE7, 8'hF2, 8'hBD},
{8'hE9, 8'hF6, 8'hC1},
{8'hE4, 8'hF1, 8'hBF},
{8'hE5, 8'hF1, 8'hC3},
{8'hD4, 8'hE0, 8'hB2},
{8'hA7, 8'hB3, 8'h82},
{8'hD5, 8'hE2, 8'hAD},
{8'hE8, 8'hF5, 8'hBE},
{8'hDE, 8'hE8, 8'hB4},
{8'h87, 8'h8F, 8'h62},
{8'h8E, 8'h93, 8'h70},
{8'hEA, 8'hEC, 8'hD5},
{8'hFD, 8'hFC, 8'hEF},
{8'hFD, 8'hFD, 8'hF1},
{8'hF9, 8'hF5, 8'hEA},
{8'hF8, 8'hF5, 8'hEA},
{8'hFD, 8'hFA, 8'hED},
{8'hF6, 8'hF5, 8'hDB},
{8'hEE, 8'hEF, 8'hCC},
{8'hEE, 8'hEE, 8'hD1},
{8'hF8, 8'hF5, 8'hE3},
{8'hF0, 8'hEC, 8'hDF},
{8'hEA, 8'hE8, 8'hD2},
{8'hDB, 8'hDA, 8'hBB},
{8'hD5, 8'hDC, 8'hB3},
{8'hE1, 8'hE8, 8'hB8},
{8'hBB, 8'hC2, 8'h8F},
{8'hBE, 8'hC2, 8'h9A},
{8'hDC, 8'hDC, 8'hC4},
{8'hF3, 8'hF1, 8'hE4},
{8'hE9, 8'hE6, 8'hD5},
{8'hEB, 8'hE9, 8'hD0},
{8'hE3, 8'hDD, 8'hC3},
{8'hE8, 8'hE3, 8'hCC},
{8'hEE, 8'hE9, 8'hD9},
{8'hF3, 8'hEE, 8'hE6},
{8'hD0, 8'hCB, 8'hCC},
{8'h38, 8'h33, 8'h3E},
{8'h1C, 8'h19, 8'h2A},
{8'h87, 8'h83, 8'h97},
{8'hD3, 8'hD0, 8'hD3},
{8'hFD, 8'hFC, 8'hFD},
{8'hFF, 8'hFF, 8'hFF},
{8'hFF, 8'hFF, 8'hFF},
{8'hFF, 8'hFF, 8'hFF},
{8'hF7, 8'hF6, 8'hF7},
{8'hF5, 8'hF4, 8'hF5},
{8'hD2, 8'hCF, 8'hD0},
{8'h98, 8'h8D, 8'h9B},
{8'h66, 8'h61, 8'h84},
{8'h25, 8'h34, 8'h75},
{8'h1E, 8'h47, 8'h9C},
{8'h19, 8'h54, 8'hAD},
{8'h13, 8'h58, 8'hB2},
{8'h0E, 8'h57, 8'hBA},
{8'h0E, 8'h56, 8'hC0},
{8'h15, 8'h55, 8'hB7},
{8'h18, 8'h4A, 8'h9D},
{8'h08, 8'h1A, 8'h56},
{8'h02, 8'h01, 8'h25},
{8'h08, 8'h02, 8'h16},
{8'h0B, 8'h06, 8'h17},
{8'h00, 8'h00, 8'h11},
{8'h3D, 8'h46, 8'h5C},
{8'hDC, 8'hDC, 8'hC4},
{8'hB2, 8'hB1, 8'h91},
{8'h8F, 8'h8E, 8'h6F},
{8'hD8, 8'hD5, 8'hC2},
{8'hCA, 8'hC6, 8'hBE},
{8'hBC, 8'hB8, 8'hB0},
{8'hD7, 8'hD5, 8'hBE},
{8'hEE, 8'hEE, 8'hCA},
{8'hE8, 8'hE6, 8'hD2},
{8'hFC, 8'hF9, 8'hDF},
{8'hDE, 8'hD8, 8'hB8},
{8'hDA, 8'hCE, 8'hB5},
{8'hFA, 8'hEE, 8'hE1},
{8'hFE, 8'hF6, 8'hEF},
{8'hED, 8'hE7, 8'hD7},
{8'hDB, 8'hDA, 8'hC2},
{8'hF7, 8'hFA, 8'hEC},
{8'hFA, 8'hFA, 8'hEB},
{8'hF4, 8'hEF, 8'hE2},
{8'hF8, 8'hEC, 8'hEC},
{8'hED, 8'hE0, 8'hE7},
{8'hED, 8'hE8, 8'hE6},
{8'hEF, 8'hF8, 8'hDC},
{8'hB4, 8'hC4, 8'h95},
{8'hB0, 8'hB5, 8'h9A},
{8'hEE, 8'hF4, 8'hCB},
{8'hEC, 8'hF4, 8'hBC},
{8'hEA, 8'hF2, 8'hBD},
{8'h8F, 8'h95, 8'h74},
{8'h76, 8'h77, 8'h70},
{8'h7C, 8'h7B, 8'h84},
{8'h7A, 8'h78, 8'h84},
{8'h7C, 8'h7B, 8'h7C},
{8'h7F, 8'h7D, 8'h7D},
{8'h7E, 8'h7C, 8'h7D},
{8'h81, 8'h7F, 8'h80},
{8'h7E, 8'h7C, 8'h7D},
{8'h7E, 8'h7C, 8'h7D},
{8'h7F, 8'h7D, 8'h7E},
{8'h7F, 8'h7D, 8'h7E},
{8'h81, 8'h7C, 8'h7F},
{8'h83, 8'h7D, 8'h80},
{8'h82, 8'h7C, 8'h7F},
{8'h81, 8'h7D, 8'h80},
{8'h7F, 8'h7D, 8'h83},
{8'h7D, 8'h7D, 8'h85},
{8'h7A, 8'h7E, 8'h89},
{8'h79, 8'h7E, 8'h89},
{8'h7F, 8'h7D, 8'h7F},
{8'h80, 8'h7C, 8'h7E},
{8'h80, 8'h7D, 8'h7E},
{8'h80, 8'h7D, 8'h7E},
{8'h80, 8'h7D, 8'h7E},
{8'h80, 8'h7D, 8'h7E},
{8'h80, 8'h7D, 8'h7E},
{8'h80, 8'h7D, 8'h7E},
{8'h7F, 8'h7D, 8'h7D},
{8'h7F, 8'h7E, 8'h7F},
{8'h7D, 8'h7E, 8'h80},
{8'h7D, 8'h7E, 8'h81},
{8'h7D, 8'h7E, 8'h81},
{8'h7E, 8'h7F, 8'h81},
{8'h7F, 8'h7F, 8'h80},
{8'h7E, 8'h7D, 8'h7A},
{8'hA5, 8'hAD, 8'h8A},
{8'hEE, 8'hFC, 8'hC0},
{8'hE1, 8'hF8, 8'hAF},
{8'hDB, 8'hF3, 8'hB8},
{8'hDF, 8'hF4, 8'hC2},
{8'hE3, 8'hF4, 8'hBA},
{8'hE7, 8'hF2, 8'hB2},
{8'hEA, 8'hF1, 8'hB5},
{8'hE6, 8'hF4, 8'hB8},
{8'hE5, 8'hF3, 8'hBA},
{8'hDE, 8'hEB, 8'hB7},
{8'hD4, 8'hE0, 8'hB0},
{8'hD4, 8'hE0, 8'hB2},
{8'hD2, 8'hDE, 8'hAF},
{8'hCA, 8'hD6, 8'hA3},
{8'hC7, 8'hD4, 8'h9F},
{8'hD5, 8'hDD, 8'hAD},
{8'hD3, 8'hD9, 8'hAE},
{8'hD7, 8'hDB, 8'hB5},
{8'hF4, 8'hF7, 8'hD8},
{8'hF7, 8'hF8, 8'hE2},
{8'hF9, 8'hF8, 8'hEA},
{8'hFB, 8'hFA, 8'hF0},
{8'hFD, 8'hFC, 8'hF5},
{8'hFF, 8'hFF, 8'hF5},
{8'hF9, 8'hF7, 8'hF4},
{8'hF4, 8'hF1, 8'hEA},
{8'hF6, 8'hF5, 8'hE3},
{8'hF9, 8'hF9, 8'hE7},
{8'hEC, 8'hE9, 8'hDF},
{8'hDA, 8'hD8, 8'hC6},
{8'hBE, 8'hBF, 8'h9D},
{8'hC7, 8'hD0, 8'hA4},
{8'hED, 8'hF6, 8'hC3},
{8'hDA, 8'hE4, 8'hAC},
{8'hB8, 8'hBF, 8'h91},
{8'hD6, 8'hD8, 8'hBE},
{8'hFB, 8'hFA, 8'hEC},
{8'hEA, 8'hE8, 8'hDA},
{8'hEF, 8'hEE, 8'hD9},
{8'hDF, 8'hDE, 8'hBF},
{8'hF0, 8'hEE, 8'hD3},
{8'hEB, 8'hEA, 8'hD7},
{8'hF2, 8'hEF, 8'hE5},
{8'hBF, 8'hBB, 8'hB9},
{8'h68, 8'h64, 8'h69},
{8'h50, 8'h4D, 8'h55},
{8'hCD, 8'hCA, 8'hD3},
{8'hFB, 8'hFA, 8'hFB},
{8'hFB, 8'hFB, 8'hFB},
{8'hFB, 8'hFA, 8'hFB},
{8'hFE, 8'hFD, 8'hFE},
{8'hFD, 8'hFC, 8'hFD},
{8'hE8, 8'hE5, 8'hE6},
{8'hFD, 8'hFC, 8'hFD},
{8'hFF, 8'hFF, 8'hFF},
{8'hF1, 8'hEA, 8'hFA},
{8'h7C, 8'h86, 8'hB4},
{8'h1D, 8'h24, 8'h5F},
{8'h3C, 8'h42, 8'h7A},
{8'h2E, 8'h4E, 8'h90},
{8'h19, 8'h50, 8'h9C},
{8'h19, 8'h58, 8'hB0},
{8'h0E, 8'h53, 8'hB8},
{8'h1E, 8'h58, 8'hB3},
{8'h12, 8'h32, 8'h79},
{8'h00, 8'h00, 8'h2B},
{8'h07, 8'h01, 8'h19},
{8'h06, 8'h01, 8'h0E},
{8'h04, 8'h04, 8'h10},
{8'h0E, 8'h11, 8'h1F},
{8'hBE, 8'hC6, 8'hCD},
{8'hBF, 8'hBE, 8'hAA},
{8'hA3, 8'hA0, 8'h87},
{8'hBF, 8'hBD, 8'hA7},
{8'hF8, 8'hF4, 8'hEA},
{8'hFE, 8'hF8, 8'hFD},
{8'hFF, 8'hF8, 8'hFE},
{8'hF9, 8'hF5, 8'hEE},
{8'hF0, 8'hEE, 8'hDA},
{8'hE9, 8'hE4, 8'hD2},
{8'hE4, 8'hE0, 8'hC7},
{8'hD2, 8'hCD, 8'hB1},
{8'hF4, 8'hEF, 8'hDB},
{8'hFE, 8'hF7, 8'hF0},
{8'hFC, 8'hF6, 8'hF2},
{8'hEA, 8'hE7, 8'hDA},
{8'hCC, 8'hCD, 8'hB6},
{8'hF2, 8'hF5, 8'hE6},
{8'hE4, 8'hE6, 8'hD2},
{8'hE6, 8'hE3, 8'hCF},
{8'hF4, 8'hEE, 8'hE3},
{8'hE9, 8'hE3, 8'hE0},
{8'hE5, 8'hE4, 8'hDD},
{8'hE2, 8'hEB, 8'hD0},
{8'h98, 8'hA8, 8'h7F},
{8'h75, 8'h78, 8'h6B},
{8'hC4, 8'hC8, 8'hAB},
{8'hF0, 8'hF7, 8'hC6},
{8'hEC, 8'hF4, 8'hC1},
{8'hA8, 8'hAD, 8'h8D},
{8'h8C, 8'h8D, 8'h86},
{8'h8C, 8'h89, 8'h92},
{8'h7C, 8'h79, 8'h86},
{8'h82, 8'h80, 8'h82},
{8'h7E, 8'h7C, 8'h7C},
{8'h7D, 8'h7B, 8'h7C},
{8'h7F, 8'h7D, 8'h7E},
{8'h7F, 8'h7D, 8'h7E},
{8'h7E, 8'h7C, 8'h7D},
{8'h7E, 8'h7C, 8'h7D},
{8'h7E, 8'h7C, 8'h7D},
{8'h88, 8'h78, 8'h85},
{8'h88, 8'h78, 8'h85},
{8'h87, 8'h77, 8'h86},
{8'h87, 8'h77, 8'h87},
{8'h87, 8'h78, 8'h87},
{8'h87, 8'h78, 8'h87},
{8'h87, 8'h78, 8'h87},
{8'h86, 8'h78, 8'h87},
{8'h83, 8'h7C, 8'h7D},
{8'h82, 8'h7C, 8'h7C},
{8'h82, 8'h7C, 8'h7C},
{8'h82, 8'h7C, 8'h7C},
{8'h82, 8'h7C, 8'h7C},
{8'h82, 8'h7C, 8'h7C},
{8'h82, 8'h7C, 8'h7C},
{8'h82, 8'h7C, 8'h7C},
{8'h7F, 8'h7D, 8'h81},
{8'hFF, 8'hD7, 8'h00},
{8'h80, 8'h7D, 8'h80},
{8'h80, 8'h7D, 8'h80},
{8'h80, 8'h7D, 8'h80},
{8'h80, 8'h7D, 8'h80},
{8'h7F, 8'h7D, 8'h81},
{8'h85, 8'h84, 8'h86},
{8'hD6, 8'hEC, 8'hCC},
{8'hE1, 8'hFC, 8'hC9},
{8'hDA, 8'hF8, 8'hB7},
{8'hDC, 8'hF8, 8'hB8},
{8'hDE, 8'hF5, 8'hBB},
{8'hE3, 8'hF3, 8'hBE},
{8'hE7, 8'hF2, 8'hB9},
{8'hE9, 8'hF1, 8'hB6},
{8'hE4, 8'hF0, 8'hB9},
{8'hE3, 8'hF0, 8'hBD},
{8'hE2, 8'hEE, 8'hC0},
{8'hE0, 8'hEC, 8'hC1},
{8'hE2, 8'hED, 8'hC3},
{8'hE7, 8'hF2, 8'hC6},
{8'hE5, 8'hF1, 8'hC2},
{8'hDD, 8'hE8, 8'hB8},
{8'hD3, 8'hD7, 8'hAD},
{8'hD3, 8'hD7, 8'hAE},
{8'hDC, 8'hE0, 8'hB6},
{8'hE1, 8'hE6, 8'hBF},
{8'hF9, 8'hFC, 8'hDC},
{8'hF2, 8'hF5, 8'hDD},
{8'hF6, 8'hF6, 8'hE8},
{8'hF9, 8'hF9, 8'hEE},
{8'hFE, 8'hFA, 8'hE9},
{8'hFD, 8'hF5, 8'hFB},
{8'hFC, 8'hF4, 8'hFD},
{8'hFB, 8'hF8, 8'hEA},
{8'hF6, 8'hF5, 8'hE0},
{8'hF3, 8'hF1, 8'hE8},
{8'hDD, 8'hDC, 8'hCF},
{8'hB7, 8'hB9, 8'h97},
{8'hA7, 8'hB0, 8'h8C},
{8'hE3, 8'hEC, 8'hBF},
{8'hEA, 8'hF4, 8'hBF},
{8'hD3, 8'hDB, 8'hAE},
{8'hEB, 8'hEE, 8'hD5},
{8'hF3, 8'hF3, 8'hE7},
{8'hF1, 8'hF0, 8'hE6},
{8'hE0, 8'hDE, 8'hCF},
{8'hE4, 8'hE7, 8'hC6},
{8'hD6, 8'hD9, 8'hBC},
{8'hED, 8'hEE, 8'hDC},
{8'hF9, 8'hF8, 8'hF2},
{8'h7A, 8'h78, 8'h7A},
{8'h37, 8'h33, 8'h3A},
{8'h5D, 8'h58, 8'h63},
{8'hD4, 8'hCF, 8'hDA},
{8'hFC, 8'hFC, 8'hFC},
{8'hFF, 8'hFF, 8'hFF},
{8'hFF, 8'hFF, 8'hFF},
{8'hFF, 8'hFF, 8'hFF},
{8'hFF, 8'hFF, 8'hFF},
{8'hE8, 8'hE4, 8'hE5},
{8'hFA, 8'hF5, 8'hF7},
{8'hFF, 8'hFF, 8'hFF},
{8'hFF, 8'hFC, 8'hFF},
{8'h65, 8'h7E, 8'hB0},
{8'h32, 8'h42, 8'h7C},
{8'h88, 8'h86, 8'hB3},
{8'h46, 8'h61, 8'h9C},
{8'h06, 8'h34, 8'h7A},
{8'h11, 8'h3A, 8'h83},
{8'h24, 8'h52, 8'hA5},
{8'h26, 8'h52, 8'hA0},
{8'h07, 8'h14, 8'h4D},
{8'h05, 8'h01, 8'h22},
{8'h07, 8'h01, 8'h11},
{8'h04, 8'h03, 8'h12},
{8'h00, 8'h01, 8'h0B},
{8'h7C, 8'h80, 8'h87},
{8'hF5, 8'hF5, 8'hF4},
{8'hDA, 8'hD7, 8'hC8},
{8'hC7, 8'hC5, 8'hAF},
{8'hD0, 8'hCE, 8'hB5},
{8'hF0, 8'hEE, 8'hDF},
{8'hFC, 8'hF7, 8'hF8},
{8'hFB, 8'hF4, 8'hFD},
{8'hF8, 8'hF2, 8'hF5},
{8'hFB, 8'hF6, 8'hF0},
{8'hF4, 8'hEC, 8'hE3},
{8'hD0, 8'hCA, 8'hB9},
{8'hEA, 8'hE6, 8'hD2},
{8'hFF, 8'hFE, 8'hF2},
{8'hFA, 8'hF7, 8'hF5},
{8'hFF, 8'hFD, 8'hFC},
{8'hE1, 8'hE2, 8'hD6},
{8'hC5, 8'hC8, 8'hB1},
{8'hF2, 8'hF2, 8'hE8},
{8'hEB, 8'hEA, 8'hD7},
{8'hE6, 8'hE5, 8'hC6},
{8'hE8, 8'hE6, 8'hC9},
{8'hDF, 8'hDC, 8'hC9},
{8'hD8, 8'hD8, 8'hC8},
{8'hDA, 8'hDF, 8'hC9},
{8'h8C, 8'h97, 8'h79},
{8'h79, 8'h79, 8'h77},
{8'h80, 8'h82, 8'h71},
{8'hCA, 8'hD0, 8'hAC},
{8'hF3, 8'hF9, 8'hD4},
{8'hCE, 8'hD1, 8'hBA},
{8'hC0, 8'hC1, 8'hBC},
{8'hEA, 8'hE9, 8'hED},
{8'hB3, 8'hB2, 8'hB6},
{8'h77, 8'h75, 8'h76},
{8'h7F, 8'h7D, 8'h7E},
{8'h7C, 8'h7A, 8'h7B},
{8'h7E, 8'h7C, 8'h7D},
{8'h84, 8'h82, 8'h83},
{8'h7F, 8'h7D, 8'h7E},
{8'h7D, 8'h7B, 8'h7C},
{8'h7F, 8'h7D, 8'h7E},
{8'h80, 8'h7C, 8'h83},
{8'h80, 8'h7C, 8'h83},
{8'h80, 8'h7C, 8'h84},
{8'h80, 8'h7C, 8'h84},
{8'h82, 8'h7B, 8'h82},
{8'h84, 8'h7B, 8'h7F},
{8'h86, 8'h7A, 8'h7B},
{8'h87, 8'h7A, 8'h7A},
{8'h81, 8'h7C, 8'h81},
{8'h80, 8'h7C, 8'h81},
{8'h80, 8'h7C, 8'h81},
{8'h80, 8'h7C, 8'h81},
{8'h80, 8'h7C, 8'h81},
{8'h80, 8'h7C, 8'h81},
{8'h80, 8'h7C, 8'h81},
{8'h80, 8'h7C, 8'h81},
{8'h80, 8'h7C, 8'h83},
{8'h81, 8'h7C, 8'h82},
{8'h83, 8'h7B, 8'h80},
{8'h83, 8'h7B, 8'h80},
{8'h83, 8'h7B, 8'h80},
{8'h83, 8'h7C, 8'h81},
{8'h81, 8'h7C, 8'h82},
{8'h84, 8'h81, 8'h87},
{8'hAE, 8'hB1, 8'hA0},
{8'hD7, 8'hDE, 8'hBF},
{8'hE0, 8'hED, 8'hBA},
{8'hE0, 8'hF1, 8'hB1},
{8'hE1, 8'hF4, 8'hBA},
{8'hE2, 8'hF2, 8'hC4},
{8'hE3, 8'hF2, 8'hC1},
{8'hE4, 8'hF4, 8'hB8},
{8'hE4, 8'hF0, 8'hC0},
{8'hDF, 8'hEA, 8'hBF},
{8'hDC, 8'hE7, 8'hBF},
{8'hDE, 8'hE9, 8'hC3},
{8'hDB, 8'hE6, 8'hC0},
{8'hDC, 8'hE8, 8'hBE},
{8'hDF, 8'hEB, 8'hBD},
{8'hE0, 8'hEC, 8'hBC},
{8'hE9, 8'hEB, 8'hC4},
{8'hDA, 8'hDC, 8'hB3},
{8'hD0, 8'hD3, 8'hA6},
{8'hD0, 8'hD4, 8'hA7},
{8'hC1, 8'hC5, 8'h9D},
{8'hD1, 8'hD5, 8'hB6},
{8'hEF, 8'hF3, 8'hDE},
{8'hF6, 8'hF8, 8'hE6},
{8'hF5, 8'hEE, 8'hD1},
{8'hFD, 8'hEF, 8'hF6},
{8'hFF, 8'hF2, 8'hFF},
{8'hFF, 8'hF9, 8'hEC},
{8'hF9, 8'hF7, 8'hDE},
{8'hF3, 8'hF1, 8'hEB},
{8'hE6, 8'hE6, 8'hDE},
{8'hDC, 8'hE1, 8'hC0},
{8'h9B, 8'hA3, 8'h89},
{8'hBD, 8'hC8, 8'hA3},
{8'hDC, 8'hE5, 8'hB7},
{8'hE3, 8'hEA, 8'hC3},
{8'hED, 8'hF1, 8'hDB},
{8'hF0, 8'hF0, 8'hE9},
{8'hD6, 8'hD6, 8'hD1},
{8'hAE, 8'hAE, 8'hA2},
{8'hBC, 8'hC1, 8'hA3},
{8'hB4, 8'hB7, 8'h9F},
{8'hF1, 8'hF2, 8'hE8},
{8'hE3, 8'hE1, 8'hE6},
{8'h21, 8'h1F, 8'h2D},
{8'h16, 8'h11, 8'h25},
{8'h89, 8'h7F, 8'h97},
{8'h8F, 8'h88, 8'h99},
{8'h79, 8'h7B, 8'h7B},
{8'h86, 8'h89, 8'h87},
{8'hAB, 8'hAC, 8'hAB},
{8'hB2, 8'hB1, 8'hB2},
{8'hA2, 8'h9F, 8'h9F},
{8'h96, 8'h91, 8'h92},
{8'h9A, 8'h92, 8'h95},
{8'hB2, 8'hAC, 8'hAB},
{8'hB6, 8'hAB, 8'hA2},
{8'h36, 8'h57, 8'h8A},
{8'h15, 8'h34, 8'h78},
{8'h52, 8'h62, 8'h97},
{8'h2B, 8'h5A, 8'hA0},
{8'h16, 8'h4F, 8'h9A},
{8'h06, 8'h17, 8'h4F},
{8'h0B, 8'h17, 8'h51},
{8'h11, 8'h2F, 8'h72},
{8'h02, 8'h09, 8'h3A},
{8'h09, 8'h03, 8'h1E},
{8'h08, 8'h02, 8'h12},
{8'h01, 8'h04, 8'h15},
{8'h29, 8'h33, 8'h41},
{8'hE6, 8'hE9, 8'hE9},
{8'hF8, 8'hEE, 8'hE2},
{8'hF3, 8'hEF, 8'hDE},
{8'hDC, 8'hDA, 8'hBF},
{8'hC5, 8'hC6, 8'hA0},
{8'hC8, 8'hC7, 8'hA7},
{8'hF7, 8'hF5, 8'hE6},
{8'hFB, 8'hF5, 8'hF5},
{8'hFA, 8'hF4, 8'hF7},
{8'hFB, 8'hF4, 8'hF4},
{8'hF8, 8'hEF, 8'hEE},
{8'hE4, 8'hDD, 8'hD6},
{8'hF6, 8'hF2, 8'hE7},
{8'hF7, 8'hF5, 8'hF1},
{8'hF5, 8'hF5, 8'hFA},
{8'hF9, 8'hFA, 8'hFC},
{8'hD6, 8'hD8, 8'hCB},
{8'hC9, 8'hCD, 8'hB5},
{8'hE9, 8'hE5, 8'hE2},
{8'hF3, 8'hF0, 8'hDC},
{8'hCD, 8'hCB, 8'hA2},
{8'hBC, 8'hBC, 8'h8B},
{8'hD7, 8'hD8, 8'hB2},
{8'hEC, 8'hED, 8'hD4},
{8'hEA, 8'hEC, 8'hD8},
{8'hE9, 8'hEC, 8'hDA},
{8'hA5, 8'hA4, 8'hAB},
{8'h87, 8'h89, 8'h82},
{8'h8E, 8'h91, 8'h7B},
{8'hCF, 8'hD3, 8'hBB},
{8'hE6, 8'hE8, 8'hDC},
{8'hCF, 8'hCF, 8'hCD},
{8'hF0, 8'hF0, 8'hEE},
{8'hDC, 8'hDE, 8'hD7},
{8'hA5, 8'hA3, 8'hA3},
{8'h90, 8'h8E, 8'h8F},
{8'h7C, 8'h7A, 8'h7B},
{8'h80, 8'h7E, 8'h7F},
{8'h81, 8'h7F, 8'h80},
{8'h7B, 8'h79, 8'h7B},
{8'h7F, 8'h7D, 8'h7E},
{8'h89, 8'h87, 8'h89},
{8'h7A, 8'h80, 8'h80},
{8'h7A, 8'h80, 8'h80},
{8'h7A, 8'h80, 8'h81},
{8'h7A, 8'h7F, 8'h80},
{8'h7C, 8'h7F, 8'h7E},
{8'h7D, 8'h7F, 8'h7C},
{8'h7F, 8'h7F, 8'h79},
{8'h81, 8'h7E, 8'h79},
{8'h7E, 8'h7D, 8'h82},
{8'h7E, 8'h7D, 8'h83},
{8'h7E, 8'h7D, 8'h83},
{8'h7E, 8'h7D, 8'h83},
{8'h7E, 8'h7D, 8'h83},
{8'h7E, 8'h7D, 8'h83},
{8'h7E, 8'h7D, 8'h83},
{8'h7E, 8'h7D, 8'h83},
{8'h80, 8'h7C, 8'h82},
{8'h80, 8'h7C, 8'h81},
{8'h82, 8'h7C, 8'h80},
{8'h83, 8'h7B, 8'h7F},
{8'h83, 8'h7B, 8'h7F},
{8'h82, 8'h7C, 8'h81},
{8'h81, 8'h7D, 8'h82},
{8'h81, 8'h7D, 8'h82},
{8'h7C, 8'h76, 8'h6F},
{8'h84, 8'h82, 8'h70},
{8'hD4, 8'hD9, 8'hB4},
{8'hEB, 8'hF5, 8'hC0},
{8'hE4, 8'hF3, 8'hBB},
{8'hE2, 8'hF2, 8'hC1},
{8'hE0, 8'hF4, 8'hBE},
{8'hE0, 8'hF5, 8'hB9},
{8'hE1, 8'hEA, 8'hC9},
{8'hDD, 8'hE3, 8'hC7},
{8'hE5, 8'hEC, 8'hD1},
{8'hED, 8'hF4, 8'hDA},
{8'hE7, 8'hEC, 8'hD3},
{8'hE8, 8'hEE, 8'hD3},
{8'hEC, 8'hF2, 8'hD7},
{8'hF1, 8'hF8, 8'hDC},
{8'hF4, 8'hF5, 8'hE1},
{8'hF4, 8'hF7, 8'hDC},
{8'hE0, 8'hE5, 8'hBD},
{8'hD0, 8'hD6, 8'hA5},
{8'hC8, 8'hCF, 8'h9F},
{8'hBE, 8'hC4, 8'h9E},
{8'hB2, 8'hB4, 8'h9D},
{8'hF1, 8'hF2, 8'hE1},
{8'hEC, 8'hE6, 8'hC4},
{8'hF5, 8'hEA, 8'hE5},
{8'hFD, 8'hF2, 8'hF6},
{8'hEF, 8'hEA, 8'hDC},
{8'hE0, 8'hDF, 8'hC6},
{8'hFA, 8'hFA, 8'hEC},
{8'hE8, 8'hE9, 8'hDF},
{8'hD6, 8'hDA, 8'hC4},
{8'hB7, 8'hBD, 8'hA6},
{8'hD0, 8'hD7, 8'hBA},
{8'hC0, 8'hC8, 8'hA2},
{8'hE4, 8'hEC, 8'hC4},
{8'hEF, 8'hF4, 8'hD2},
{8'hD4, 8'hD7, 8'hC0},
{8'h9C, 8'h9D, 8'h8F},
{8'h91, 8'h91, 8'h86},
{8'hB8, 8'hBC, 8'hA9},
{8'hEA, 8'hEB, 8'hE2},
{8'hFD, 8'hFC, 8'hF7},
{8'h8F, 8'h8B, 8'h9B},
{8'h00, 8'h00, 8'h07},
{8'h2A, 8'h23, 8'h3F},
{8'h93, 8'h8E, 8'hA2},
{8'h9E, 8'h9B, 8'hAA},
{8'h9D, 8'h9F, 8'h9F},
{8'hAE, 8'hB0, 8'hAE},
{8'hC3, 8'hC5, 8'hC5},
{8'hA2, 8'hA2, 8'hA2},
{8'h6C, 8'h6A, 8'h6D},
{8'h65, 8'h5F, 8'h65},
{8'h86, 8'h7D, 8'h86},
{8'hCA, 8'hC0, 8'hC4},
{8'hBE, 8'hC0, 8'hBD},
{8'h15, 8'h45, 8'h7F},
{8'h0A, 8'h3C, 8'h8A},
{8'h1C, 8'h4F, 8'hA3},
{8'h11, 8'h55, 8'hB6},
{8'h19, 8'h53, 8'hA7},
{8'h21, 8'h3F, 8'h80},
{8'h06, 8'h0C, 8'h3D},
{8'h00, 8'h0B, 8'h3A},
{8'h0E, 8'h15, 8'h38},
{8'h08, 8'h01, 8'h16},
{8'h08, 8'h02, 8'h14},
{8'h06, 8'h06, 8'h1B},
{8'hAB, 8'hB4, 8'hC2},
{8'hFC, 8'hFF, 8'hFC},
{8'hFD, 8'hF5, 8'hE4},
{8'hF5, 8'hF3, 8'hDC},
{8'hD1, 8'hD2, 8'hB5},
{8'hB7, 8'hB8, 8'h95},
{8'hAF, 8'hB0, 8'h91},
{8'hC9, 8'hC8, 8'hB4},
{8'hFD, 8'hFB, 8'hF2},
{8'hF3, 8'hEF, 8'hEA},
{8'hF3, 8'hEF, 8'hEA},
{8'hF8, 8'hEB, 8'hEE},
{8'hF1, 8'hE7, 8'hE0},
{8'hF7, 8'hF2, 8'hE2},
{8'hF9, 8'hF7, 8'hE8},
{8'hF3, 8'hF3, 8'hED},
{8'hEF, 8'hF0, 8'hED},
{8'hDD, 8'hE0, 8'hD6},
{8'hE2, 8'hE6, 8'hD2},
{8'hEC, 8'hE7, 8'hE2},
{8'hD7, 8'hD3, 8'hBE},
{8'hCB, 8'hC8, 8'hA0},
{8'hE6, 8'hE4, 8'hB5},
{8'hEF, 8'hEE, 8'hC6},
{8'hE8, 8'hE6, 8'hCE},
{8'hF5, 8'hF4, 8'hE7},
{8'hFA, 8'hF9, 8'hF1},
{8'hF5, 8'hF2, 8'hF6},
{8'hE7, 8'hE5, 8'hE2},
{8'hEE, 8'hEE, 8'hE1},
{8'hF2, 8'hF3, 8'hE5},
{8'hFA, 8'hFB, 8'hF4},
{8'hF6, 8'hF6, 8'hF5},
{8'hEF, 8'hEF, 8'hEE},
{8'hD0, 8'hD1, 8'hCC},
{8'hEB, 8'hEA, 8'hE9},
{8'hAF, 8'hAD, 8'hAE},
{8'h7C, 8'h7A, 8'h7D},
{8'h82, 8'h80, 8'h83},
{8'h7E, 8'h7C, 8'h7F},
{8'h78, 8'h76, 8'h76},
{8'h87, 8'h86, 8'h82},
{8'h90, 8'h8F, 8'h89},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'h7C, 8'h7E, 8'h7D},
{8'h7B, 8'h80, 8'h76},
{8'hC8, 8'hD1, 8'hB9},
{8'hE9, 8'hF5, 8'hCE},
{8'hE1, 8'hF0, 8'hBD},
{8'hE1, 8'hF3, 8'hB8},
{8'hE2, 8'hF4, 8'hB7},
{8'hE0, 8'hF2, 8'hB8},
{8'hE6, 8'hEA, 8'hD9},
{8'hE8, 8'hEA, 8'hDE},
{8'hDD, 8'hDE, 8'hD3},
{8'hF3, 8'hF2, 8'hEA},
{8'hFC, 8'hFA, 8'hF4},
{8'hFF, 8'hFE, 8'hFA},
{8'hFF, 8'hFD, 8'hFA},
{8'hFC, 8'hF9, 8'hF5},
{8'hF8, 8'hFA, 8'hF7},
{8'hF3, 8'hF7, 8'hE9},
{8'hE0, 8'hE7, 8'hC6},
{8'hDC, 8'hE4, 8'hB6},
{8'hD7, 8'hDF, 8'hAE},
{8'hB0, 8'hB6, 8'h8E},
{8'h97, 8'h99, 8'h80},
{8'hC6, 8'hC7, 8'hB6},
{8'hDF, 8'hDE, 8'hC0},
{8'hE5, 8'hE4, 8'hCD},
{8'hEF, 8'hED, 8'hDF},
{8'hC4, 8'hC3, 8'hB3},
{8'hD0, 8'hD2, 8'hB9},
{8'hDE, 8'hE2, 8'hC4},
{8'hE1, 8'hE4, 8'hCF},
{8'hDF, 8'hE1, 8'hD6},
{8'hD2, 8'hD5, 8'hBF},
{8'hDC, 8'hDF, 8'hCA},
{8'hE6, 8'hE9, 8'hD4},
{8'hBF, 8'hC5, 8'hA3},
{8'hAF, 8'hB7, 8'h88},
{8'hC6, 8'hCD, 8'hA1},
{8'h9A, 8'h9E, 8'h84},
{8'hAE, 8'hB0, 8'hA6},
{8'hF4, 8'hF5, 8'hED},
{8'hFB, 8'hF9, 8'hF9},
{8'hE8, 8'hE5, 8'hE4},
{8'h49, 8'h42, 8'h56},
{8'h2A, 8'h27, 8'h2E},
{8'h5E, 8'h5B, 8'h6E},
{8'hD5, 8'hD6, 8'hD9},
{8'hFA, 8'hFD, 8'hFC},
{8'hFF, 8'hFF, 8'hFF},
{8'hFF, 8'hFF, 8'hFF},
{8'hFF, 8'hFF, 8'hFF},
{8'hFF, 8'hFF, 8'hFF},
{8'hFF, 8'hFF, 8'hFF},
{8'hD4, 8'hCE, 8'hDA},
{8'hA1, 8'h94, 8'hA4},
{8'h9B, 8'h8C, 8'h9D},
{8'h81, 8'h9B, 8'hB9},
{8'h12, 8'h45, 8'h83},
{8'h20, 8'h4E, 8'h98},
{8'h0E, 8'h56, 8'hC4},
{8'h0E, 8'h56, 8'hCA},
{8'h20, 8'h4F, 8'hAC},
{8'h1F, 8'h56, 8'hB4},
{8'h15, 8'h33, 8'h75},
{8'h00, 8'h03, 8'h21},
{8'h05, 8'h06, 8'h1F},
{8'h09, 8'h01, 8'h15},
{8'h05, 8'h00, 8'h0F},
{8'h67, 8'h65, 8'h78},
{8'hF3, 8'hF5, 8'hFF},
{8'hED, 8'hEF, 8'hED},
{8'hF7, 8'hF7, 8'hE8},
{8'hEF, 8'hF1, 8'hD6},
{8'hC6, 8'hC8, 8'hB1},
{8'hA1, 8'hA3, 8'h93},
{8'hCD, 8'hCD, 8'hC2},
{8'hEA, 8'hEA, 8'hE1},
{8'hF4, 8'hF4, 8'hE9},
{8'hF3, 8'hF3, 8'hE6},
{8'hF5, 8'hF4, 8'hE6},
{8'hFA, 8'hEE, 8'hDF},
{8'hF4, 8'hEA, 8'hCC},
{8'hF9, 8'hF4, 8'hC7},
{8'hF2, 8'hF0, 8'hC3},
{8'hF2, 8'hF1, 8'hD5},
{8'hEA, 8'hEB, 8'hDF},
{8'hF4, 8'hF6, 8'hF1},
{8'hF8, 8'hFB, 8'hF4},
{8'hF6, 8'hF4, 8'hEB},
{8'hEC, 8'hE8, 8'hD9},
{8'hED, 8'hE9, 8'hD0},
{8'hEC, 8'hE6, 8'hC9},
{8'hEA, 8'hE4, 8'hC5},
{8'hC3, 8'hBE, 8'hA6},
{8'hD6, 8'hD2, 8'hC5},
{8'hFB, 8'hF7, 8'hF1},
{8'hFC, 8'hF7, 8'hF2},
{8'hFF, 8'hFB, 8'hF5},
{8'hFF, 8'hFD, 8'hF4},
{8'hFF, 8'hFE, 8'hF4},
{8'hFF, 8'hFF, 8'hF7},
{8'hFB, 8'hFB, 8'hF7},
{8'hF1, 8'hF1, 8'hF4},
{8'hE9, 8'hE8, 8'hEE},
{8'hE9, 8'hE7, 8'hEA},
{8'hB1, 8'hAF, 8'hB0},
{8'h75, 8'h74, 8'h73},
{8'h7C, 8'h7B, 8'h77},
{8'h79, 8'h78, 8'h72},
{8'h8A, 8'h89, 8'h82},
{8'h9A, 8'h9A, 8'h92},
{8'h7A, 8'h7A, 8'h72},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'h7D, 8'h7D, 8'h81},
{8'h79, 8'h7C, 8'h77},
{8'hAB, 8'hB2, 8'hA0},
{8'hE8, 8'hF2, 8'hD1},
{8'hE1, 8'hEE, 8'hC1},
{8'hE1, 8'hF1, 8'hBA},
{8'hE1, 8'hF3, 8'hB7},
{8'hE2, 8'hF4, 8'hB9},
{8'hEA, 8'hEF, 8'hD5},
{8'hE2, 8'hE4, 8'hD3},
{8'hE7, 8'hE8, 8'hE0},
{8'hF0, 8'hEF, 8'hEE},
{8'hF0, 8'hEF, 8'hEF},
{8'hF1, 8'hEE, 8'hEB},
{8'hEA, 8'hE6, 8'hDD},
{8'hE0, 8'hDD, 8'hCE},
{8'hE2, 8'hE2, 8'hD1},
{8'hE7, 8'hE8, 8'hD1},
{8'hE8, 8'hEB, 8'hCD},
{8'hDC, 8'hE2, 8'hBD},
{8'hD3, 8'hDA, 8'hB3},
{8'hC1, 8'hC8, 8'hA4},
{8'hA3, 8'hAB, 8'h8A},
{8'hD4, 8'hDB, 8'hBD},
{8'hEB, 8'hEB, 8'hD7},
{8'hEF, 8'hED, 8'hE2},
{8'hD9, 8'hD9, 8'hD2},
{8'hA3, 8'hA5, 8'h96},
{8'hC3, 8'hC9, 8'hA9},
{8'hE6, 8'hEE, 8'hC5},
{8'hDF, 8'hE7, 8'hC4},
{8'hD0, 8'hD7, 8'hBC},
{8'hBA, 8'hBD, 8'hAA},
{8'hDB, 8'hDD, 8'hD3},
{8'hF0, 8'hF0, 8'hEC},
{8'hF1, 8'hF3, 8'hEA},
{8'hE0, 8'hE2, 8'hCF},
{8'hE5, 8'hE9, 8'hD1},
{8'hD3, 8'hD5, 8'hC7},
{8'hF7, 8'hF7, 8'hF4},
{8'hFB, 8'hFC, 8'hF3},
{8'hFC, 8'hFD, 8'hF6},
{8'h81, 8'h7D, 8'h8A},
{8'h52, 8'h50, 8'h55},
{8'h4D, 8'h48, 8'h61},
{8'hC5, 8'hC4, 8'hC9},
{8'hFF, 8'hFF, 8'hFF},
{8'hF9, 8'hFA, 8'hFA},
{8'hFE, 8'hFF, 8'hFD},
{8'hFE, 8'hFF, 8'hFF},
{8'hFC, 8'hFF, 8'hFF},
{8'hFE, 8'hFF, 8'hFF},
{8'hFF, 8'hFF, 8'hFF},
{8'hED, 8'hE4, 8'hEB},
{8'hDE, 8'hCC, 8'hD7},
{8'hF1, 8'hDB, 8'hE7},
{8'h8B, 8'h91, 8'hA4},
{8'h10, 8'h29, 8'h59},
{8'h3E, 8'h53, 8'h8B},
{8'h28, 8'h59, 8'hB3},
{8'h19, 8'h54, 8'hBB},
{8'h21, 8'h51, 8'hAE},
{8'h0F, 8'h53, 8'hBB},
{8'h1C, 8'h51, 8'hA6},
{8'h0F, 8'h20, 8'h52},
{8'h00, 8'h00, 8'h23},
{8'h02, 8'h00, 8'h12},
{8'h15, 8'h0F, 8'h19},
{8'hD7, 8'hD5, 8'hDE},
{8'hF7, 8'hFA, 8'hFF},
{8'hF0, 8'hF1, 8'hF1},
{8'hEA, 8'hE7, 8'hDF},
{8'hD3, 8'hD4, 8'hC1},
{8'hC6, 8'hC7, 8'hB7},
{8'hD9, 8'hD9, 8'hCE},
{8'hF4, 8'hF4, 8'hED},
{8'hF7, 8'hF6, 8'hF1},
{8'hFC, 8'hFB, 8'hF6},
{8'hF5, 8'hF5, 8'hEE},
{8'hEE, 8'hED, 8'hE0},
{8'hFB, 8'hF4, 8'hC0},
{8'hEB, 8'hE6, 8'hA3},
{8'hE5, 8'hE2, 8'h9B},
{8'hE7, 8'hE5, 8'hA9},
{8'hF3, 8'hF1, 8'hCE},
{8'hF0, 8'hED, 8'hE2},
{8'hF8, 8'hF5, 8'hF6},
{8'hF7, 8'hF4, 8'hF7},
{8'hF6, 8'hF3, 8'hF9},
{8'hF3, 8'hF0, 8'hF1},
{8'hEC, 8'hEA, 8'hE1},
{8'hE9, 8'hE7, 8'hD2},
{8'hEA, 8'hE7, 8'hCB},
{8'hE8, 8'hE5, 8'hC8},
{8'hEB, 8'hE9, 8'hCB},
{8'hF6, 8'hF5, 8'hDA},
{8'hFD, 8'hF9, 8'hEF},
{8'hFC, 8'hF8, 8'hEF},
{8'hF9, 8'hF5, 8'hEC},
{8'hF5, 8'hF4, 8'hEB},
{8'hF7, 8'hF7, 8'hEF},
{8'hFE, 8'hFF, 8'hFA},
{8'hFF, 8'hFF, 8'hFD},
{8'hF5, 8'hF6, 8'hF6},
{8'hDE, 8'hDC, 8'hE5},
{8'hA0, 8'h9F, 8'h9D},
{8'hA3, 8'hA4, 8'h8F},
{8'hC3, 8'hC7, 8'hA5},
{8'hBA, 8'hBD, 8'h9D},
{8'h9E, 8'h9F, 8'h8E},
{8'h80, 8'h7E, 8'h82},
{8'h7E, 8'h79, 8'h8C},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'h7F, 8'h7D, 8'h81},
{8'h7A, 8'h79, 8'h83},
{8'h82, 8'h83, 8'h85},
{8'h7C, 8'h80, 8'h76},
{8'hB8, 8'hC0, 8'hA8},
{8'hE6, 8'hF1, 8'hCB},
{8'hE5, 8'hF3, 8'hC3},
{8'hE2, 8'hF3, 8'hBA},
{8'hE1, 8'hF2, 8'hB9},
{8'hE1, 8'hE8, 8'hC4},
{8'hDD, 8'hE0, 8'hCA},
{8'hEE, 8'hEF, 8'hE7},
{8'hFB, 8'hF9, 8'hFD},
{8'hF9, 8'hF6, 8'hF9},
{8'hF7, 8'hF3, 8'hF2},
{8'hEE, 8'hEA, 8'hDC},
{8'hE1, 8'hDF, 8'hC7},
{8'hDF, 8'hDB, 8'hC2},
{8'hF7, 8'hF5, 8'hE0},
{8'hFD, 8'hFD, 8'hEA},
{8'hF5, 8'hF6, 8'hE5},
{8'hDF, 8'hE2, 8'hD0},
{8'hD8, 8'hE1, 8'hC8},
{8'h97, 8'hA4, 8'h84},
{8'hBC, 8'hCA, 8'hA7},
{8'hF7, 8'hF8, 8'hEF},
{8'hF5, 8'hF4, 8'hF3},
{8'hC2, 8'hC2, 8'hC1},
{8'h89, 8'h8D, 8'h7D},
{8'hBC, 8'hC4, 8'h9D},
{8'hE3, 8'hF0, 8'hBB},
{8'hEA, 8'hF8, 8'hC2},
{8'hD2, 8'hDF, 8'hB1},
{8'hC7, 8'hCB, 8'hB3},
{8'hF6, 8'hF7, 8'hF0},
{8'hFF, 8'hFE, 8'hFF},
{8'hFC, 8'hF9, 8'hFF},
{8'hFE, 8'hFE, 8'hFD},
{8'hF8, 8'hF9, 8'hEE},
{8'hF2, 8'hF4, 8'hE8},
{8'hF7, 8'hF7, 8'hF2},
{8'hFC, 8'hFD, 8'hF5},
{8'hBE, 8'hC1, 8'hB9},
{8'h11, 8'h10, 8'h23},
{8'h25, 8'h27, 8'h29},
{8'h5E, 8'h5C, 8'h7A},
{8'hEF, 8'hF0, 8'hEF},
{8'hF4, 8'hF2, 8'hF5},
{8'hFE, 8'hFD, 8'hF7},
{8'hFD, 8'hFF, 8'hFD},
{8'hFC, 8'hFF, 8'hFF},
{8'hFD, 8'hFF, 8'hFF},
{8'hFF, 8'hFF, 8'hFF},
{8'hFF, 8'hFD, 8'hFE},
{8'hF0, 8'hE4, 8'hE8},
{8'hE4, 8'hCD, 8'hD3},
{8'hE9, 8'hCE, 8'hD7},
{8'h7F, 8'h86, 8'hA2},
{8'h28, 8'h42, 8'h74},
{8'h85, 8'h91, 8'hC2},
{8'h32, 8'h56, 8'hA5},
{8'h20, 8'h52, 8'hAF},
{8'h1D, 8'h4E, 8'hAA},
{8'h03, 8'h52, 8'hC3},
{8'h0E, 8'h56, 8'hBC},
{8'h1E, 8'h3E, 8'h87},
{8'h01, 8'h08, 8'h3B},
{8'h01, 8'h02, 8'h18},
{8'h1A, 8'h16, 8'h1A},
{8'hDC, 8'hDB, 8'hDA},
{8'hF2, 8'hF5, 8'hF5},
{8'hF6, 8'hF7, 8'hF7},
{8'hEC, 8'hE8, 8'hE6},
{8'hD9, 8'hD9, 8'hCC},
{8'hF5, 8'hF6, 8'hEB},
{8'hFE, 8'hFD, 8'hF8},
{8'hF5, 8'hF4, 8'hF3},
{8'hFA, 8'hF9, 8'hF8},
{8'hFB, 8'hFA, 8'hF8},
{8'hF7, 8'hF6, 8'hF2},
{8'hF1, 8'hF0, 8'hE4},
{8'hFA, 8'hF5, 8'hB2},
{8'hE0, 8'hDB, 8'h8B},
{8'hD4, 8'hD2, 8'h81},
{8'hE8, 8'hE6, 8'hA5},
{8'hF5, 8'hF0, 8'hCC},
{8'hF7, 8'hEF, 8'hE5},
{8'hFE, 8'hF8, 8'hF8},
{8'hF9, 8'hF3, 8'hF6},
{8'hF7, 8'hF5, 8'hFD},
{8'hEF, 8'hEF, 8'hF3},
{8'hEF, 8'hF0, 8'hED},
{8'hE7, 8'hE9, 8'hDC},
{8'hEC, 8'hEE, 8'hD8},
{8'hDE, 8'hDE, 8'hC0},
{8'hE8, 8'hE7, 8'hC2},
{8'hF0, 8'hEE, 8'hC7},
{8'hF6, 8'hF2, 8'hE2},
{8'hF5, 8'hF2, 8'hE5},
{8'hF5, 8'hF2, 8'hE8},
{8'hF3, 8'hF2, 8'hEA},
{8'hEE, 8'hEE, 8'hE6},
{8'hF4, 8'hF5, 8'hEC},
{8'hF6, 8'hF7, 8'hED},
{8'hF3, 8'hF5, 8'hEA},
{8'hF4, 8'hF3, 8'hF1},
{8'hE8, 8'hE8, 8'hDA},
{8'hEF, 8'hF3, 8'hD0},
{8'hF4, 8'hFA, 8'hCB},
{8'hBC, 8'hC1, 8'h98},
{8'h78, 8'h79, 8'h66},
{8'h82, 8'h7F, 8'h88},
{8'h7F, 8'h79, 8'h94},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'h80, 8'h7E, 8'h82},
{8'h82, 8'h7F, 8'h8B},
{8'h7D, 8'h7B, 8'h82},
{8'h7E, 8'h7F, 8'h7D},
{8'h7E, 8'h82, 8'h73},
{8'hC6, 8'hCE, 8'hB3},
{8'hBF, 8'hCA, 8'hA3},
{8'hDC, 8'hE9, 8'hBA},
{8'hE5, 8'hF2, 8'hC0},
{8'hE4, 8'hEB, 8'hC2},
{8'hE6, 8'hEB, 8'hCE},
{8'hF1, 8'hF3, 8'hE7},
{8'hF6, 8'hF4, 8'hF6},
{8'hF6, 8'hF3, 8'hF6},
{8'hF2, 8'hEE, 8'hE8},
{8'hE5, 8'hE3, 8'hCE},
{8'hE1, 8'hDF, 8'hC0},
{8'hEA, 8'hE4, 8'hCF},
{8'hFF, 8'hFB, 8'hEF},
{8'hFA, 8'hF3, 8'hF2},
{8'hFB, 8'hF8, 8'hFB},
{8'hFA, 8'hFC, 8'hFE},
{8'hE4, 8'hEB, 8'hE6},
{8'hC2, 8'hCF, 8'hBC},
{8'hCA, 8'hD8, 8'hBE},
{8'hF7, 8'hF8, 8'hF7},
{8'hF6, 8'hF5, 8'hFB},
{8'hCC, 8'hCD, 8'hCE},
{8'h8E, 8'h92, 8'h82},
{8'hCB, 8'hD6, 8'hAB},
{8'hE1, 8'hF0, 8'hB1},
{8'hE5, 8'hF4, 8'hB4},
{8'hD2, 8'hE1, 8'hA6},
{8'hC2, 8'hC6, 8'hA2},
{8'hED, 8'hEE, 8'hDF},
{8'hFE, 8'hFC, 8'hFE},
{8'hFA, 8'hF7, 8'hFD},
{8'hFA, 8'hF9, 8'hF7},
{8'hF9, 8'hF9, 8'hEB},
{8'hF9, 8'hFA, 8'hE7},
{8'hF2, 8'hF4, 8'hE3},
{8'hE0, 8'hE1, 8'hDE},
{8'h37, 8'h37, 8'h3C},
{8'h00, 8'h00, 8'h0E},
{8'h06, 8'h08, 8'h1B},
{8'h9F, 8'hA1, 8'hB4},
{8'hEA, 8'hEB, 8'hF3},
{8'hEC, 8'hE9, 8'hEC},
{8'hFE, 8'hFD, 8'hF7},
{8'hFD, 8'hFF, 8'hFE},
{8'hFC, 8'hFF, 8'hFF},
{8'hFD, 8'hFF, 8'hFF},
{8'hFF, 8'hFE, 8'hFF},
{8'hFC, 8'hF9, 8'hFA},
{8'hFB, 8'hF0, 8'hF4},
{8'hE5, 8'hCD, 8'hD2},
{8'hDC, 8'hC3, 8'hCD},
{8'h4B, 8'h6C, 8'hA6},
{8'h1C, 8'h4E, 8'h98},
{8'h5A, 8'h76, 8'hB5},
{8'h28, 8'h53, 8'hA6},
{8'h1D, 8'h51, 8'hAD},
{8'h1D, 8'h4E, 8'hA9},
{8'h06, 8'h5A, 8'hCD},
{8'h0B, 8'h58, 8'hC5},
{8'h22, 8'h4E, 8'hAA},
{8'h0D, 8'h21, 8'h63},
{8'h00, 8'h01, 8'h1E},
{8'h07, 8'h06, 8'h08},
{8'hC0, 8'hC0, 8'hBA},
{8'hF7, 8'hFA, 8'hF5},
{8'hF1, 8'hF1, 8'hEE},
{8'hF4, 8'hF0, 8'hEE},
{8'hEF, 8'hEE, 8'hE5},
{8'hFB, 8'hFB, 8'hF4},
{8'hF9, 8'hF8, 8'hF5},
{8'hFE, 8'hFD, 8'hFC},
{8'hF3, 8'hF2, 8'hF1},
{8'hFB, 8'hFB, 8'hF8},
{8'hF6, 8'hF5, 8'hEF},
{8'hF1, 8'hF0, 8'hE5},
{8'hF9, 8'hF2, 8'hC6},
{8'hE6, 8'hDF, 8'hA8},
{8'hDE, 8'hD9, 8'h9F},
{8'hF3, 8'hED, 8'hBE},
{8'hF6, 8'hEE, 8'hD5},
{8'hF9, 8'hF0, 8'hE8},
{8'hFA, 8'hF1, 8'hEE},
{8'hF6, 8'hEF, 8'hE9},
{8'hBE, 8'hC0, 8'hB2},
{8'hA7, 8'hA9, 8'h9E},
{8'hB8, 8'hBC, 8'hB3},
{8'hE5, 8'hE9, 8'hE0},
{8'hF0, 8'hF2, 8'hE4},
{8'hE4, 8'hE2, 8'hCB},
{8'hEC, 8'hE8, 8'hC6},
{8'hF6, 8'hF0, 8'hCA},
{8'hF5, 8'hF3, 8'hDB},
{8'hF8, 8'hF5, 8'hE3},
{8'hFB, 8'hF9, 8'hEE},
{8'hFD, 8'hFB, 8'hF6},
{8'hF5, 8'hF4, 8'hF0},
{8'hEE, 8'hEF, 8'hE4},
{8'hEB, 8'hEE, 8'hDB},
{8'hE7, 8'hEC, 8'hD3},
{8'hEE, 8'hF2, 8'hD1},
{8'hEB, 8'hEF, 8'hCC},
{8'hF0, 8'hF5, 8'hD1},
{8'hE9, 8'hEC, 8'hCC},
{8'h8D, 8'h8F, 8'h78},
{8'h78, 8'h78, 8'h6E},
{8'h7D, 8'h7B, 8'h7D},
{8'h7D, 8'h7B, 8'h84},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'h7F, 8'h7D, 8'h81},
{8'h7F, 8'h7C, 8'h85},
{8'h7F, 8'h7C, 8'h84},
{8'h7E, 8'h7E, 8'h80},
{8'h7D, 8'h7E, 8'h79},
{8'h84, 8'h88, 8'h79},
{8'h83, 8'h8A, 8'h70},
{8'h9F, 8'hA9, 8'h87},
{8'hDC, 8'hE7, 8'hBF},
{8'hE8, 8'hF0, 8'hC5},
{8'hF2, 8'hF7, 8'hD4},
{8'hF3, 8'hF6, 8'hE0},
{8'hEA, 8'hEB, 8'hDE},
{8'hF2, 8'hF1, 8'hE6},
{8'hE4, 8'hE3, 8'hD1},
{8'hDC, 8'hDB, 8'hBF},
{8'hD7, 8'hD6, 8'hB5},
{8'hE5, 8'hDF, 8'hD1},
{8'hFE, 8'hFA, 8'hF6},
{8'hFB, 8'hF5, 8'hFB},
{8'hFD, 8'hF9, 8'hFF},
{8'hF8, 8'hF7, 8'hFF},
{8'hF1, 8'hF6, 8'hF7},
{8'hB1, 8'hBA, 8'hB4},
{8'hEC, 8'hF5, 8'hE9},
{8'hF4, 8'hF2, 8'hF2},
{8'hFA, 8'hF7, 8'hFC},
{8'hEF, 8'hED, 8'hED},
{8'hB7, 8'hB9, 8'hA7},
{8'hC6, 8'hCE, 8'hA0},
{8'hD7, 8'hE3, 8'hA2},
{8'hE8, 8'hF6, 8'hB2},
{8'hD3, 8'hE0, 8'hA1},
{8'hD1, 8'hD4, 8'hAA},
{8'hE7, 8'hE7, 8'hCF},
{8'hF5, 8'hF3, 8'hEC},
{8'hFB, 8'hF9, 8'hF4},
{8'hF9, 8'hF8, 8'hE8},
{8'hF9, 8'hFA, 8'hE0},
{8'hF4, 8'hF4, 8'hD8},
{8'hF4, 8'hF5, 8'hDC},
{8'h57, 8'h58, 8'h5D},
{8'h00, 8'h00, 8'h13},
{8'h00, 8'h04, 8'h13},
{8'h1D, 8'h22, 8'h4E},
{8'hC7, 8'hCE, 8'hDE},
{8'hD4, 8'hD3, 8'hF0},
{8'hF7, 8'hF5, 8'hF2},
{8'hFE, 8'hF9, 8'hF4},
{8'hFE, 8'hFE, 8'hFF},
{8'hFE, 8'hFF, 8'hFF},
{8'hFD, 8'hFF, 8'hFF},
{8'hFE, 8'hFF, 8'hFF},
{8'hFD, 8'hFB, 8'hFD},
{8'hFE, 8'hF7, 8'hFD},
{8'hEB, 8'hD8, 8'hE2},
{8'hCD, 8'hBC, 8'hCD},
{8'h1F, 8'h5E, 8'hB4},
{8'h0A, 8'h58, 8'hBD},
{8'h1B, 8'h4C, 8'hA0},
{8'h18, 8'h54, 8'hB2},
{8'h15, 8'h52, 8'hB3},
{8'h1D, 8'h50, 8'hAA},
{8'h07, 8'h56, 8'hC5},
{8'h0F, 8'h54, 8'hBD},
{8'h1B, 8'h50, 8'hB7},
{8'h16, 8'h37, 8'h84},
{8'h00, 8'h01, 8'h28},
{8'h01, 8'h01, 8'h06},
{8'h97, 8'h97, 8'h92},
{8'hF8, 8'hFB, 8'hF3},
{8'hF7, 8'hF7, 8'hEE},
{8'hEB, 8'hE7, 8'hDD},
{8'hD2, 8'hD2, 8'hC6},
{8'hFE, 8'hFE, 8'hF4},
{8'hFC, 8'hFC, 8'hF6},
{8'hF8, 8'hF7, 8'hF2},
{8'hF6, 8'hF6, 8'hF0},
{8'hFA, 8'hFA, 8'hF1},
{8'hED, 8'hEE, 8'hDF},
{8'hF1, 8'hF2, 8'hE2},
{8'hF8, 8'hF0, 8'hE8},
{8'hF7, 8'hF0, 8'hDF},
{8'hEE, 8'hE8, 8'hCE},
{8'hFB, 8'hF5, 8'hDE},
{8'hFB, 8'hF3, 8'hE9},
{8'hF7, 8'hEE, 8'hEA},
{8'hF9, 8'hF1, 8'hE8},
{8'hF6, 8'hF1, 8'hDD},
{8'hB3, 8'hB7, 8'h8F},
{8'h96, 8'h9C, 8'h7B},
{8'h7C, 8'h83, 8'h6E},
{8'h88, 8'h8E, 8'h81},
{8'hE1, 8'hE3, 8'hD5},
{8'hE6, 8'hE3, 8'hCB},
{8'hF5, 8'hEC, 8'hC5},
{8'hFC, 8'hF0, 8'hC2},
{8'hF3, 8'hF2, 8'hD3},
{8'hF7, 8'hF5, 8'hDF},
{8'hFC, 8'hF9, 8'hEE},
{8'hFE, 8'hFC, 8'hF9},
{8'hFA, 8'hF9, 8'hF5},
{8'hF4, 8'hF6, 8'hE8},
{8'hEA, 8'hEE, 8'hD2},
{8'hCD, 8'hD5, 8'hAD},
{8'hE7, 8'hF0, 8'hB2},
{8'hEA, 8'hF1, 8'hBE},
{8'hF5, 8'hF8, 8'hDC},
{8'hBC, 8'hBC, 8'hB2},
{8'h7C, 8'h7B, 8'h7B},
{8'h80, 8'h7F, 8'h7E},
{8'h7F, 8'h7F, 8'h77},
{8'h7D, 8'h7D, 8'h70},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'h81, 8'h7C, 8'h80},
{8'h7F, 8'h7D, 8'h81},
{8'h7F, 8'h7D, 8'h82},
{8'h7F, 8'h7E, 8'h80},
{8'h81, 8'h81, 8'h7F},
{8'h7E, 8'h81, 8'h76},
{8'h89, 8'h8F, 8'h7B},
{8'hA4, 8'hAD, 8'h92},
{8'hD1, 8'hD9, 8'hB1},
{8'hDD, 8'hE3, 8'hBB},
{8'hDB, 8'hE2, 8'hBC},
{8'hD7, 8'hDB, 8'hB7},
{8'hE6, 8'hE9, 8'hC8},
{8'hE1, 8'hE2, 8'hC1},
{8'hDC, 8'hDC, 8'hBD},
{8'hCD, 8'hCC, 8'hAE},
{8'hD2, 8'hD1, 8'hC1},
{8'hF5, 8'hF4, 8'hEA},
{8'hF7, 8'hF5, 8'hF0},
{8'hF9, 8'hF9, 8'hF9},
{8'hFC, 8'hFC, 8'hFB},
{8'hFE, 8'hFF, 8'hFD},
{8'hC7, 8'hCB, 8'hC6},
{8'hEF, 8'hF2, 8'hEC},
{8'hF9, 8'hF3, 8'hEC},
{8'hFB, 8'hF4, 8'hF2},
{8'hF7, 8'hF1, 8'hED},
{8'hBD, 8'hBB, 8'hA6},
{8'hCC, 8'hCF, 8'hA2},
{8'hD4, 8'hDB, 8'h9E},
{8'hE2, 8'hEB, 8'hAC},
{8'hD9, 8'hE1, 8'hA7},
{8'hCB, 8'hCC, 8'hA9},
{8'hDE, 8'hDC, 8'hC6},
{8'hED, 8'hEB, 8'hDC},
{8'hF8, 8'hF6, 8'hE5},
{8'hFA, 8'hF9, 8'hDE},
{8'hFD, 8'hFE, 8'hE0},
{8'hF0, 8'hEF, 8'hD5},
{8'h81, 8'h7F, 8'h70},
{8'h00, 8'h00, 8'h0E},
{8'h04, 8'h07, 8'h25},
{8'h05, 8'h0B, 8'h26},
{8'h13, 8'h18, 8'h4D},
{8'h84, 8'h8B, 8'hA7},
{8'hD4, 8'hD2, 8'hF4},
{8'hFB, 8'hF5, 8'hF4},
{8'hFF, 8'hFA, 8'hF7},
{8'hFF, 8'hFE, 8'hFD},
{8'hFF, 8'hFF, 8'hFD},
{8'hFD, 8'hFF, 8'hFF},
{8'hFB, 8'hFF, 8'hFF},
{8'hFA, 8'hFD, 8'hFF},
{8'hFF, 8'hFF, 8'hFF},
{8'hE1, 8'hD8, 8'hE8},
{8'h84, 8'h7C, 8'h95},
{8'h0B, 8'h4A, 8'hA7},
{8'h07, 8'h56, 8'hC3},
{8'h17, 8'h50, 8'hAB},
{8'h10, 8'h55, 8'hBB},
{8'h11, 8'h55, 8'hBA},
{8'h1C, 8'h50, 8'hAB},
{8'h0B, 8'h55, 8'hC0},
{8'h15, 8'h52, 8'hB6},
{8'h11, 8'h51, 8'hBA},
{8'h1B, 8'h46, 8'h99},
{8'h02, 8'h05, 8'h36},
{8'h00, 8'h00, 8'h13},
{8'h34, 8'h32, 8'h37},
{8'hE6, 8'hE8, 8'hE1},
{8'hF5, 8'hF6, 8'hE5},
{8'hF0, 8'hED, 8'hD5},
{8'hEE, 8'hEF, 8'hDB},
{8'hF6, 8'hF7, 8'hE6},
{8'hF1, 8'hF2, 8'hE4},
{8'hEC, 8'hED, 8'hDF},
{8'hF0, 8'hF1, 8'hE2},
{8'hF3, 8'hF4, 8'hE1},
{8'hD1, 8'hD3, 8'hB9},
{8'hBB, 8'hBE, 8'hA4},
{8'hDA, 8'hD5, 8'hDB},
{8'hFC, 8'hF9, 8'hF6},
{8'hF4, 8'hF2, 8'hE6},
{8'hF5, 8'hF1, 8'hE8},
{8'hFC, 8'hF7, 8'hF6},
{8'hF9, 8'hF4, 8'hF5},
{8'hFB, 8'hF6, 8'hF0},
{8'hF2, 8'hEF, 8'hDB},
{8'hA2, 8'hA2, 8'h75},
{8'hAA, 8'hAC, 8'h88},
{8'h86, 8'h89, 8'h74},
{8'h9D, 8'hA1, 8'h92},
{8'hE5, 8'hE6, 8'hD1},
{8'hF5, 8'hF0, 8'hC7},
{8'hF2, 8'hE5, 8'hA4},
{8'hF8, 8'hEB, 8'h9E},
{8'hF2, 8'hF1, 8'hCA},
{8'hF4, 8'hF2, 8'hD9},
{8'hF9, 8'hF6, 8'hEB},
{8'hFD, 8'hFA, 8'hF8},
{8'hF4, 8'hF3, 8'hEF},
{8'hF2, 8'hF5, 8'hE3},
{8'hEB, 8'hF1, 8'hCD},
{8'hC9, 8'hD2, 8'hA0},
{8'hE8, 8'hF0, 8'hB3},
{8'hE9, 8'hEF, 8'hBE},
{8'hB8, 8'hBB, 8'hA0},
{8'h7C, 8'h7C, 8'h74},
{8'h7E, 8'h7C, 8'h7D},
{8'h7E, 8'h7D, 8'h7D},
{8'h7D, 8'h7C, 8'h76},
{8'h7E, 8'h7E, 8'h71},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'h81, 8'h7D, 8'h7A},
{8'h81, 8'h7D, 8'h7D},
{8'h7F, 8'h7D, 8'h81},
{8'h7E, 8'h7C, 8'h83},
{8'h7D, 8'h7D, 8'h82},
{8'h7F, 8'h81, 8'h7F},
{8'h7D, 8'h80, 8'h77},
{8'h7A, 8'h7E, 8'h70},
{8'hAB, 8'hB2, 8'h8E},
{8'hD1, 8'hD8, 8'hAB},
{8'hCA, 8'hD3, 8'h9D},
{8'hD8, 8'hE1, 8'hA7},
{8'hD8, 8'hDD, 8'hA6},
{8'hD5, 8'hD8, 8'hAA},
{8'hCF, 8'hCE, 8'hAD},
{8'hB4, 8'hB3, 8'h9A},
{8'hB6, 8'hBC, 8'hA2},
{8'hE1, 8'hE6, 8'hCB},
{8'hF0, 8'hF4, 8'hD9},
{8'hEC, 8'hF0, 8'hD5},
{8'hEB, 8'hEF, 8'hD6},
{8'hF7, 8'hFA, 8'hE7},
{8'hE3, 8'hE5, 8'hD7},
{8'hEC, 8'hEC, 8'hE1},
{8'hF8, 8'hEF, 8'hDF},
{8'hFB, 8'hF1, 8'hE8},
{8'hFB, 8'hF3, 8'hEA},
{8'hE2, 8'hDC, 8'hC4},
{8'hD1, 8'hD0, 8'hA3},
{8'hD2, 8'hD4, 8'h9A},
{8'hDD, 8'hE0, 8'hA7},
{8'hDE, 8'hE1, 8'hB1},
{8'hE4, 8'hE1, 8'hD0},
{8'hF8, 8'hF5, 8'hEA},
{8'hF8, 8'hF5, 8'hE9},
{8'hF1, 8'hEE, 8'hD9},
{8'hF2, 8'hF2, 8'hD3},
{8'hFF, 8'hFF, 8'hE4},
{8'hA7, 8'hA4, 8'h94},
{8'h0D, 8'h07, 8'h0A},
{8'h04, 8'h04, 8'h1D},
{8'h04, 8'h05, 8'h24},
{8'h0A, 8'h0F, 8'h3F},
{8'h05, 8'h0E, 8'h3D},
{8'h3C, 8'h42, 8'h74},
{8'hC3, 8'hC2, 8'hDA},
{8'hFF, 8'hF6, 8'hFE},
{8'hFF, 8'hF9, 8'hF8},
{8'hFF, 8'hFE, 8'hF9},
{8'hFF, 8'hFF, 8'hFC},
{8'hFF, 8'hFF, 8'hFF},
{8'hFF, 8'hFF, 8'hFF},
{8'hF3, 8'hF9, 8'hFB},
{8'hB5, 8'hB9, 8'hC6},
{8'h3C, 8'h3C, 8'h54},
{8'h07, 8'h07, 8'h25},
{8'h1F, 8'h45, 8'h96},
{8'h10, 8'h4E, 8'hAE},
{8'h16, 8'h45, 8'h99},
{8'h10, 8'h56, 8'hBB},
{8'h0D, 8'h56, 8'hBD},
{8'h1A, 8'h51, 8'hAC},
{8'h0C, 8'h54, 8'hBF},
{8'h18, 8'h51, 8'hB4},
{8'h0F, 8'h56, 8'hBE},
{8'h19, 8'h4B, 8'hA1},
{8'h05, 8'h11, 8'h4B},
{8'h02, 8'h00, 8'h23},
{8'h02, 8'h01, 8'h0D},
{8'h90, 8'h91, 8'h8B},
{8'hEC, 8'hED, 8'hD3},
{8'hED, 8'hED, 8'hC8},
{8'hED, 8'hEF, 8'hD4},
{8'hF1, 8'hF4, 8'hDA},
{8'hEB, 8'hED, 8'hD5},
{8'hF0, 8'hF2, 8'hDA},
{8'hE0, 8'hE3, 8'hC8},
{8'hC3, 8'hC7, 8'hA7},
{8'hC3, 8'hC7, 8'hA2},
{8'hA5, 8'hAA, 8'h84},
{8'hCF, 8'hD1, 8'hC7},
{8'hFA, 8'hFE, 8'hEF},
{8'hF7, 8'hFA, 8'hE7},
{8'hF9, 8'hFA, 8'hF0},
{8'hF7, 8'hF5, 8'hF9},
{8'hFB, 8'hF8, 8'hFF},
{8'hF3, 8'hEF, 8'hF2},
{8'hF8, 8'hF6, 8'hEC},
{8'hC6, 8'hC1, 8'hA4},
{8'hB9, 8'hB5, 8'h9F},
{8'hC4, 8'hC4, 8'hB7},
{8'hF5, 8'hF8, 8'hEA},
{8'hFD, 8'hFD, 8'hDC},
{8'hF0, 8'hEA, 8'hA6},
{8'hE0, 8'hD2, 8'h67},
{8'hEC, 8'hDC, 8'h61},
{8'hF6, 8'hF5, 8'hC5},
{8'hF7, 8'hF7, 8'hDB},
{8'hFD, 8'hFA, 8'hEF},
{8'hFE, 8'hFC, 8'hFD},
{8'hF6, 8'hF6, 8'hF4},
{8'hF0, 8'hF3, 8'hE0},
{8'hE6, 8'hEE, 8'hC4},
{8'hC1, 8'hCB, 8'h94},
{8'hD8, 8'hDD, 8'hB7},
{8'h94, 8'h98, 8'h75},
{8'h92, 8'h96, 8'h75},
{8'h9B, 8'h9E, 8'h82},
{8'h96, 8'h97, 8'h83},
{8'h90, 8'h90, 8'h87},
{8'h88, 8'h86, 8'h88},
{8'h84, 8'h81, 8'h89},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'h7F, 8'h7D, 8'h7F},
{8'h7E, 8'h7C, 8'h7B},
{8'h82, 8'h7F, 8'h80},
{8'h81, 8'h7E, 8'h82},
{8'h7E, 8'h7C, 8'h81},
{8'h7E, 8'h7D, 8'h81},
{8'h7E, 8'h7E, 8'h7F},
{8'h82, 8'h83, 8'h7F},
{8'h7C, 8'h7D, 8'h77},
{8'h82, 8'h84, 8'h7A},
{8'h9E, 8'hA1, 8'h8C},
{8'h9B, 8'hA2, 8'h7B},
{8'hC6, 8'hCE, 8'h99},
{8'hE8, 8'hF0, 8'hB7},
{8'hE6, 8'hEC, 8'hB8},
{8'hE4, 8'hE7, 8'hBF},
{8'hCA, 8'hCC, 8'hAE},
{8'hCE, 8'hD2, 8'hBF},
{8'hE9, 8'hED, 8'hD9},
{8'hE2, 8'hE9, 8'hCF},
{8'hF4, 8'hFA, 8'hE1},
{8'hF0, 8'hF4, 8'hDF},
{8'hF0, 8'hF0, 8'hDE},
{8'hF2, 8'hEF, 8'hD9},
{8'hF7, 8'hF1, 8'hD6},
{8'hF5, 8'hEC, 8'hD6},
{8'hFA, 8'hF1, 8'hE3},
{8'hFB, 8'hF4, 8'hEB},
{8'hF9, 8'hF2, 8'hE4},
{8'hF2, 8'hF0, 8'hD6},
{8'hD5, 8'hD3, 8'hAD},
{8'hD3, 8'hD4, 8'hA8},
{8'hDD, 8'hDF, 8'hB4},
{8'hF4, 8'hF1, 8'hE3},
{8'hF8, 8'hF5, 8'hED},
{8'hF8, 8'hF5, 8'hE9},
{8'hEC, 8'hEC, 8'hD1},
{8'hF0, 8'hF1, 8'hCA},
{8'hD9, 8'hD9, 8'hBB},
{8'h2C, 8'h27, 8'h28},
{8'h02, 8'h00, 8'h13},
{8'h08, 8'h05, 8'h15},
{8'h04, 8'h0C, 8'h27},
{8'h09, 8'h13, 8'h41},
{8'h06, 8'h0A, 8'h2F},
{8'h21, 8'h2F, 8'h72},
{8'h63, 8'h76, 8'hA2},
{8'hEA, 8'hED, 8'hFC},
{8'hFF, 8'hFC, 8'hF8},
{8'hFF, 8'hFF, 8'hF1},
{8'hFE, 8'hFF, 8'hFF},
{8'hE2, 8'hF9, 8'hFB},
{8'hA8, 8'hC4, 8'hD7},
{8'h62, 8'h73, 8'h9F},
{8'h0E, 8'h10, 8'h3A},
{8'h00, 8'h00, 8'h18},
{8'h08, 8'h08, 8'h2C},
{8'h1E, 8'h47, 8'h84},
{8'h1E, 8'h4E, 8'hA8},
{8'h0D, 8'h30, 8'h8A},
{8'h0E, 8'h41, 8'h9E},
{8'h19, 8'h55, 8'hB7},
{8'h16, 8'h4E, 8'hB8},
{8'h0F, 8'h57, 8'hC5},
{8'h10, 8'h55, 8'hAE},
{8'h0F, 8'h55, 8'hBC},
{8'h18, 8'h4C, 8'hA5},
{8'h0D, 8'h1F, 8'h59},
{8'h00, 8'h01, 8'h1F},
{8'h00, 8'h00, 8'h0F},
{8'h2F, 8'h2B, 8'h35},
{8'hD7, 8'hD7, 8'hBE},
{8'hDD, 8'hE2, 8'hA5},
{8'hE2, 8'hE5, 8'hBE},
{8'hF4, 8'hF5, 8'hD8},
{8'hFC, 8'hFC, 8'hE8},
{8'hFF, 8'hFC, 8'hF0},
{8'hEB, 8'hEB, 8'hDC},
{8'hDC, 8'hDC, 8'hC6},
{8'hC4, 8'hC6, 8'hA6},
{8'hAA, 8'hAD, 8'h88},
{8'hDF, 8'hE2, 8'hD6},
{8'hF8, 8'hFA, 8'hEE},
{8'hF6, 8'hF8, 8'hEA},
{8'hF9, 8'hFB, 8'hF1},
{8'hF0, 8'hEF, 8'hEC},
{8'hD5, 8'hD4, 8'hD4},
{8'hF3, 8'hF2, 8'hEE},
{8'hF1, 8'hF0, 8'hE5},
{8'hF4, 8'hF0, 8'hDB},
{8'hC2, 8'hBC, 8'hAC},
{8'hDB, 8'hD8, 8'hCC},
{8'hF8, 8'hF6, 8'hE7},
{8'hFA, 8'hF8, 8'hD8},
{8'hEA, 8'hE6, 8'hAB},
{8'hD9, 8'hD1, 8'h79},
{8'hE6, 8'hDD, 8'h79},
{8'hF6, 8'hF8, 8'hCE},
{8'hFA, 8'hFB, 8'hDF},
{8'hFE, 8'hFD, 8'hEF},
{8'hFE, 8'hFD, 8'hF7},
{8'hFC, 8'hFA, 8'hF1},
{8'hFC, 8'hFC, 8'hE7},
{8'hEE, 8'hF2, 8'hC9},
{8'hB1, 8'hB6, 8'h84},
{8'hD8, 8'hDB, 8'hBF},
{8'hC1, 8'hC4, 8'hA9},
{8'hD4, 8'hD7, 8'hBA},
{8'hD2, 8'hD5, 8'hBA},
{8'h82, 8'h83, 8'h6F},
{8'h81, 8'h81, 8'h79},
{8'h81, 8'h7F, 8'h84},
{8'h80, 8'h7D, 8'h89},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'h7E, 8'h7C, 8'h80},
{8'h7F, 8'h7D, 8'h82},
{8'h81, 8'h7F, 8'h83},
{8'h7E, 8'h7C, 8'h7F},
{8'h81, 8'h7F, 8'h81},
{8'h82, 8'h80, 8'h80},
{8'h7C, 8'h7B, 8'h79},
{8'h7B, 8'h7A, 8'h77},
{8'h81, 8'h80, 8'h7E},
{8'h7D, 8'h7B, 8'h89},
{8'h77, 8'h77, 8'h7B},
{8'h82, 8'h85, 8'h76},
{8'hD3, 8'hD9, 8'hB8},
{8'hCD, 8'hD4, 8'hAA},
{8'hDE, 8'hE5, 8'hBB},
{8'hEE, 8'hF4, 8'hCF},
{8'hFA, 8'hFC, 8'hE1},
{8'hFE, 8'hFA, 8'hF7},
{8'hF9, 8'hF8, 8'hF1},
{8'hF9, 8'hFB, 8'hF4},
{8'hFC, 8'hFF, 8'hFC},
{8'hF8, 8'hF8, 8'hF9},
{8'hF3, 8'hEE, 8'hE5},
{8'hF3, 8'hEB, 8'hC9},
{8'hF8, 8'hEE, 8'hB8},
{8'hF4, 8'hEE, 8'hD0},
{8'hF7, 8'hF2, 8'hDD},
{8'hFB, 8'hF6, 8'hEB},
{8'hFA, 8'hF5, 8'hF1},
{8'hF8, 8'hF5, 8'hF0},
{8'hF4, 8'hF4, 8'hE4},
{8'hD6, 8'hD9, 8'hBB},
{8'hD4, 8'hD8, 8'hB1},
{8'hEE, 8'hEE, 8'hD7},
{8'hF3, 8'hF1, 8'hE3},
{8'hF5, 8'hF3, 8'hE4},
{8'hF0, 8'hF1, 8'hD0},
{8'hEB, 8'hEE, 8'hC2},
{8'h8E, 8'h8F, 8'h73},
{8'h02, 8'h00, 8'h0A},
{8'h0A, 8'h02, 8'h2C},
{8'h07, 8'h02, 8'h0A},
{8'h00, 8'h14, 8'h37},
{8'h04, 8'h12, 8'h33},
{8'h04, 8'h01, 8'h25},
{8'h1C, 8'h3B, 8'h87},
{8'h22, 8'h4F, 8'hA3},
{8'h8B, 8'hA2, 8'hC6},
{8'hF7, 8'hFF, 8'hFF},
{8'hE1, 8'hE6, 8'hDF},
{8'h88, 8'hA3, 8'hC8},
{8'h30, 8'h6D, 8'h9D},
{8'h17, 8'h56, 8'h8E},
{8'h1E, 8'h3B, 8'h91},
{8'h02, 8'h02, 8'h3E},
{8'h03, 8'h00, 8'h14},
{8'h05, 8'h06, 8'h2E},
{8'h0D, 8'h47, 8'h88},
{8'h20, 8'h54, 8'hB0},
{8'h18, 8'h40, 8'hA3},
{8'h03, 8'h20, 8'h6E},
{8'h17, 8'h3C, 8'h8D},
{8'h1D, 8'h4D, 8'hBA},
{8'h0F, 8'h4E, 8'hBB},
{8'h08, 8'h58, 8'hAE},
{8'h10, 8'h52, 8'hB9},
{8'h1D, 8'h50, 8'hAE},
{8'h0D, 8'h25, 8'h5D},
{8'h00, 8'h03, 8'h18},
{8'h07, 8'h03, 8'h1C},
{8'h05, 8'h00, 8'h1A},
{8'h83, 8'h82, 8'h71},
{8'hDD, 8'hE7, 8'h97},
{8'hE0, 8'hE3, 8'hB2},
{8'hF6, 8'hF5, 8'hD7},
{8'hFE, 8'hFA, 8'hEE},
{8'hFF, 8'hFC, 8'hFD},
{8'hFF, 8'hFD, 8'hFF},
{8'hFB, 8'hF7, 8'hF3},
{8'hEB, 8'hE8, 8'hD7},
{8'hC0, 8'hBF, 8'hA5},
{8'hEB, 8'hE9, 8'hE8},
{8'hF6, 8'hF4, 8'hF4},
{8'hF8, 8'hF7, 8'hF4},
{8'hFF, 8'hFF, 8'hF9},
{8'hD7, 8'hD7, 8'hCB},
{8'hA0, 8'hA1, 8'h91},
{8'hDD, 8'hDE, 8'hCB},
{8'hEE, 8'hEE, 8'hDA},
{8'hF1, 8'hED, 8'hD2},
{8'hD4, 8'hCF, 8'hB7},
{8'hD0, 8'hCB, 8'hB6},
{8'hEB, 8'hE6, 8'hD2},
{8'hED, 8'hE9, 8'hD3},
{8'hEE, 8'hEA, 8'hCE},
{8'hEA, 8'hE8, 8'hC5},
{8'hE6, 8'hE5, 8'hBE},
{8'hED, 8'hF0, 8'hD0},
{8'hF1, 8'hF5, 8'hDB},
{8'hF8, 8'hF8, 8'hE5},
{8'hFD, 8'hFA, 8'hEC},
{8'hF5, 8'hF1, 8'hE3},
{8'hF4, 8'hF0, 8'hDE},
{8'hF2, 8'hEE, 8'hD3},
{8'hC0, 8'hBC, 8'h9C},
{8'hC8, 8'hCB, 8'hAA},
{8'hE1, 8'hE3, 8'hC8},
{8'hFD, 8'hFD, 8'hED},
{8'hC1, 8'hC1, 8'hB8},
{8'h7B, 8'h79, 8'h78},
{8'h7E, 8'h7C, 8'h7E},
{8'h7D, 8'h7B, 8'h7E},
{8'h7F, 8'h7E, 8'h7F},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'h81, 8'h7F, 8'h84},
{8'h7E, 8'h7C, 8'h80},
{8'h82, 8'h80, 8'h83},
{8'hBA, 8'hB8, 8'hBA},
{8'h7E, 8'h7C, 8'h7C},
{8'hA3, 8'hA2, 8'hA0},
{8'h90, 8'h8F, 8'h8C},
{8'h74, 8'h73, 8'h70},
{8'h7E, 8'h7E, 8'h7B},
{8'h79, 8'h7A, 8'h70},
{8'h8E, 8'h92, 8'h7D},
{8'hE1, 8'hE5, 8'hC8},
{8'hE6, 8'hEB, 8'hCD},
{8'hEB, 8'hEF, 8'hD5},
{8'hF8, 8'hFA, 8'hE9},
{8'hED, 8'hEE, 8'hE3},
{8'hEF, 8'hEC, 8'hDD},
{8'hF9, 8'hF8, 8'hE8},
{8'hFD, 8'hFD, 8'hF2},
{8'hFC, 8'hFC, 8'hF6},
{8'hFC, 8'hF9, 8'hF3},
{8'hFC, 8'hF8, 8'hDF},
{8'hF9, 8'hF3, 8'hB7},
{8'hF0, 8'hEA, 8'h98},
{8'hE6, 8'hE4, 8'hB5},
{8'hF5, 8'hF2, 8'hCF},
{8'hF7, 8'hF4, 8'hDE},
{8'hF8, 8'hF5, 8'hEA},
{8'hF7, 8'hF5, 8'hED},
{8'hF6, 8'hF4, 8'hE6},
{8'hED, 8'hF0, 8'hD6},
{8'hD7, 8'hDB, 8'hBA},
{8'hDE, 8'hE0, 8'hCA},
{8'hE0, 8'hE1, 8'hD2},
{8'hDA, 8'hDB, 8'hCC},
{8'hE5, 8'hE8, 8'hCE},
{8'hE5, 8'hE8, 8'hC7},
{8'h3A, 8'h3A, 8'h2D},
{8'h00, 8'h00, 8'h0A},
{8'h09, 8'h01, 8'h2B},
{8'h07, 8'h01, 8'h1F},
{8'h08, 8'h20, 8'h55},
{8'h02, 8'h0F, 8'h3A},
{8'h01, 8'h00, 8'h26},
{8'h12, 8'h35, 8'h86},
{8'h1C, 8'h51, 8'hB3},
{8'h30, 8'h52, 8'h98},
{8'h6B, 8'h84, 8'hB1},
{8'h37, 8'h5B, 8'h8A},
{8'h17, 8'h49, 8'hA7},
{8'h13, 8'h56, 8'hB9},
{8'h19, 8'h56, 8'hA5},
{8'h10, 8'h2B, 8'h70},
{8'h00, 8'h02, 8'h24},
{8'h00, 8'h03, 8'h13},
{8'h0A, 8'h18, 8'h49},
{8'h14, 8'h44, 8'hA3},
{8'h18, 8'h50, 8'hAF},
{8'h1C, 8'h54, 8'hAC},
{8'h0D, 8'h34, 8'h7C},
{8'h00, 8'h0B, 8'h49},
{8'h17, 8'h33, 8'h78},
{8'h27, 8'h55, 8'hAE},
{8'h15, 8'h52, 8'hBD},
{8'h11, 8'h52, 8'hBB},
{8'h1D, 8'h51, 8'hB1},
{8'h0D, 8'h25, 8'h64},
{8'h00, 8'h04, 8'h21},
{8'h05, 8'h03, 8'h1F},
{8'h07, 8'h00, 8'h20},
{8'h24, 8'h21, 8'h1D},
{8'hC6, 8'hCD, 8'h8D},
{8'hED, 8'hF0, 8'hBE},
{8'hFA, 8'hFA, 8'hD7},
{8'hFC, 8'hF9, 8'hE6},
{8'hFB, 8'hF7, 8'hF2},
{8'hFC, 8'hF7, 8'hF5},
{8'hFA, 8'hF6, 8'hF0},
{8'hF3, 8'hF0, 8'hE0},
{8'hE6, 8'hE3, 8'hCE},
{8'hEE, 8'hED, 8'hE7},
{8'hF0, 8'hEF, 8'hEB},
{8'hF3, 8'hF3, 8'hEB},
{8'hF8, 8'hF8, 8'hED},
{8'hDE, 8'hDE, 8'hD1},
{8'hD1, 8'hD2, 8'hC1},
{8'hBB, 8'hBD, 8'hA9},
{8'hC9, 8'hCA, 8'hB4},
{8'hD9, 8'hD7, 8'hB7},
{8'hC4, 8'hC1, 8'hA3},
{8'hB5, 8'hB1, 8'h97},
{8'hA9, 8'hA4, 8'h8D},
{8'hA9, 8'hA5, 8'h8E},
{8'hEB, 8'hE7, 8'hCC},
{8'hE9, 8'hE6, 8'hC5},
{8'hF0, 8'hEE, 8'hCB},
{8'hEE, 8'hF0, 8'hD2},
{8'hF1, 8'hF3, 8'hDB},
{8'hF9, 8'hF8, 8'hEA},
{8'hFE, 8'hFB, 8'hF4},
{8'hFD, 8'hFA, 8'hF5},
{8'hF0, 8'hEA, 8'hE2},
{8'hE6, 8'hE0, 8'hD1},
{8'hD8, 8'hD4, 8'hBF},
{8'hED, 8'hEF, 8'hD2},
{8'hFD, 8'hFE, 8'hE6},
{8'hFD, 8'hFD, 8'hEE},
{8'hA5, 8'hA5, 8'h9D},
{8'h78, 8'h77, 8'h75},
{8'h7C, 8'h7A, 8'h7B},
{8'h82, 8'h80, 8'h81},
{8'h7F, 8'h7D, 8'h7E},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'h7E, 8'h7C, 8'h7F},
{8'h7E, 8'h7C, 8'h81},
{8'h7E, 8'h7C, 8'h80},
{8'h87, 8'h85, 8'h88},
{8'hDE, 8'hDC, 8'hDE},
{8'hA2, 8'hA1, 8'hA0},
{8'hEE, 8'hED, 8'hEB},
{8'hCB, 8'hCA, 8'hC7},
{8'hB6, 8'hB5, 8'hB1},
{8'h8E, 8'h8F, 8'h89},
{8'h8A, 8'h8B, 8'h81},
{8'hB6, 8'hB9, 8'hA9},
{8'hEE, 8'hF1, 8'hDE},
{8'hF9, 8'hFC, 8'hE9},
{8'hFC, 8'hFE, 8'hEF},
{8'hF4, 8'hF6, 8'hEA},
{8'hE3, 8'hE4, 8'hDA},
{8'hF1, 8'hEF, 8'hD5},
{8'hF5, 8'hF4, 8'hDB},
{8'hF8, 8'hF6, 8'hE5},
{8'hFA, 8'hF6, 8'hED},
{8'hFC, 8'hF6, 8'hEA},
{8'hFD, 8'hF8, 8'hD0},
{8'hED, 8'hE9, 8'h95},
{8'hD4, 8'hD3, 8'h62},
{8'hE3, 8'hE5, 8'hA4},
{8'hFD, 8'hFD, 8'hCE},
{8'hF7, 8'hF7, 8'hD6},
{8'hF1, 8'hEF, 8'hDE},
{8'hF0, 8'hEE, 8'hE3},
{8'hF4, 8'hF5, 8'hE8},
{8'hE5, 8'hE8, 8'hD4},
{8'hD5, 8'hD9, 8'hC0},
{8'hEE, 8'hF0, 8'hDA},
{8'hDE, 8'hE0, 8'hCD},
{8'hD6, 8'hD7, 8'hC7},
{8'hE4, 8'hE6, 8'hD4},
{8'hAE, 8'hB0, 8'hA0},
{8'h09, 8'h08, 8'h08},
{8'h04, 8'h01, 8'h17},
{8'h08, 8'h01, 8'h2A},
{8'h04, 8'h00, 8'h2F},
{8'h13, 8'h2D, 8'h6F},
{8'h04, 8'h11, 8'h3C},
{8'h00, 8'h00, 8'h21},
{8'h0E, 8'h37, 8'h86},
{8'h11, 8'h52, 8'hBF},
{8'h1B, 8'h4E, 8'hAF},
{8'h1B, 8'h4A, 8'h9F},
{8'h13, 8'h54, 8'hAA},
{8'h0C, 8'h52, 8'hD3},
{8'h09, 8'h4E, 8'hD6},
{8'h1C, 8'h51, 8'hB3},
{8'h0C, 8'h1D, 8'h50},
{8'h00, 8'h02, 8'h0F},
{8'h00, 8'h0A, 8'h20},
{8'h14, 8'h33, 8'h79},
{8'h1B, 8'h43, 8'hB0},
{8'h13, 8'h4F, 8'hAC},
{8'h13, 8'h58, 8'hAD},
{8'h23, 8'h57, 8'hAB},
{8'h0F, 8'h1E, 8'h5C},
{8'h00, 8'h03, 8'h28},
{8'h14, 8'h2B, 8'h68},
{8'h22, 8'h4C, 8'hB5},
{8'h19, 8'h55, 8'hB9},
{8'h20, 8'h51, 8'hB2},
{8'h0E, 8'h24, 8'h6B},
{8'h00, 8'h05, 8'h2A},
{8'h03, 8'h04, 8'h22},
{8'h07, 8'h02, 8'h26},
{8'h01, 8'h00, 8'h06},
{8'h73, 8'h78, 8'h4F},
{8'hEF, 8'hF1, 8'hC0},
{8'hFB, 8'hFB, 8'hD6},
{8'hFE, 8'hFC, 8'hE3},
{8'hFE, 8'hFC, 8'hF0},
{8'hFC, 8'hF8, 8'hF2},
{8'hF7, 8'hF2, 8'hEB},
{8'hF3, 8'hF0, 8'hE4},
{8'hDB, 8'hD8, 8'hC9},
{8'hE0, 8'hDF, 8'hD6},
{8'hEB, 8'hEB, 8'hE2},
{8'hF0, 8'hF0, 8'hE5},
{8'hE3, 8'hE3, 8'hD6},
{8'hD1, 8'hD2, 8'hC2},
{8'hD2, 8'hD3, 8'hC1},
{8'h8F, 8'h91, 8'h7D},
{8'h87, 8'h89, 8'h72},
{8'hB2, 8'hB3, 8'h8E},
{8'hB1, 8'hB1, 8'h8D},
{8'hB2, 8'hB1, 8'h91},
{8'h9F, 8'h9D, 8'h83},
{8'hA9, 8'hA7, 8'h8F},
{8'hE9, 8'hE7, 8'hD0},
{8'hF0, 8'hEE, 8'hD5},
{8'hF5, 8'hF3, 8'hDB},
{8'hF5, 8'hF7, 8'hE2},
{8'hF5, 8'hF7, 8'hE7},
{8'hF7, 8'hF6, 8'hEC},
{8'hFA, 8'hF7, 8'hF1},
{8'hFB, 8'hF7, 8'hF0},
{8'hF1, 8'hEC, 8'hDD},
{8'hD6, 8'hD1, 8'hB8},
{8'hE9, 8'hE6, 8'hC7},
{8'hFB, 8'hFD, 8'hE2},
{8'hF6, 8'hF8, 8'hE3},
{8'hEE, 8'hEF, 8'hE1},
{8'hC6, 8'hC5, 8'hBE},
{8'h82, 8'h81, 8'h80},
{8'h7F, 8'h7D, 8'h7E},
{8'h90, 8'h8E, 8'h8F},
{8'h8B, 8'h89, 8'h8A},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'h7E, 8'h7C, 8'h81},
{8'h7F, 8'h7D, 8'h81},
{8'h7D, 8'h7B, 8'h7E},
{8'hC3, 8'hC1, 8'hC4},
{8'hF9, 8'hF8, 8'hF7},
{8'hF7, 8'hF6, 8'hF4},
{8'hF9, 8'hF8, 8'hF5},
{8'hFD, 8'hFC, 8'hF8},
{8'hEC, 8'hEB, 8'hEC},
{8'hF2, 8'hF1, 8'hF2},
{8'hFD, 8'hFD, 8'hFB},
{8'hF8, 8'hF8, 8'hF1},
{8'hF6, 8'hF7, 8'hEA},
{8'hFB, 8'hFD, 8'hEB},
{8'hE4, 8'hE8, 8'hD1},
{8'hCF, 8'hD3, 8'hB8},
{8'hF3, 8'hF5, 8'hD5},
{8'hF9, 8'hFA, 8'hDD},
{8'hFC, 8'hF9, 8'hE6},
{8'hFB, 8'hF4, 8'hEA},
{8'hFE, 8'hF7, 8'hE9},
{8'hFA, 8'hF5, 8'hC8},
{8'hE1, 8'hE0, 8'h83},
{8'hC2, 8'hC5, 8'h4A},
{8'hD6, 8'hDB, 8'h92},
{8'hF3, 8'hF7, 8'hC0},
{8'hE5, 8'hE7, 8'hC1},
{8'hE5, 8'hE5, 8'hD0},
{8'hE9, 8'hEA, 8'hDE},
{8'hD9, 8'hDA, 8'hCF},
{8'hD3, 8'hD7, 8'hC5},
{8'hE5, 8'hE9, 8'hD3},
{8'hF8, 8'hFC, 8'hE1},
{8'hE0, 8'hE5, 8'hCB},
{8'hE0, 8'hE2, 8'hCE},
{8'hEA, 8'hEB, 8'hE0},
{8'h5A, 8'h5A, 8'h5B},
{8'h00, 8'h00, 8'h09},
{8'h09, 8'h06, 8'h22},
{8'h05, 8'h02, 8'h24},
{8'h07, 8'h08, 8'h40},
{8'h1D, 8'h3E, 8'h83},
{8'h03, 8'h14, 8'h39},
{8'h02, 8'h03, 8'h19},
{8'h08, 8'h36, 8'h7B},
{8'h0E, 8'h58, 8'hC3},
{8'h10, 8'h50, 8'hBA},
{8'h15, 8'h54, 8'hB9},
{8'h0B, 8'h59, 8'hB6},
{8'h07, 8'h54, 8'hD1},
{8'h0F, 8'h50, 8'hDB},
{8'h21, 8'h47, 8'hAD},
{8'h0A, 8'h16, 8'h3A},
{8'h00, 8'h01, 8'h0B},
{8'h02, 8'h0E, 8'h3D},
{8'h20, 8'h43, 8'hA3},
{8'h1A, 8'h44, 8'hA7},
{8'h0F, 8'h4F, 8'hA1},
{8'h0E, 8'h59, 8'hB6},
{8'h19, 8'h4F, 8'hC1},
{8'h2A, 8'h41, 8'h98},
{8'h06, 8'h0A, 8'h2C},
{8'h00, 8'h00, 8'h22},
{8'h0C, 8'h1C, 8'h67},
{8'h17, 8'h48, 8'h9D},
{8'h26, 8'h4D, 8'hAA},
{8'h10, 8'h24, 8'h6E},
{8'h00, 8'h03, 8'h2A},
{8'h01, 8'h01, 8'h21},
{8'h05, 8'h01, 8'h29},
{8'h03, 8'h00, 8'h12},
{8'h1E, 8'h21, 8'h12},
{8'hD5, 8'hD7, 8'hAF},
{8'hFA, 8'hFA, 8'hD7},
{8'hF9, 8'hF8, 8'hDE},
{8'hF9, 8'hF6, 8'hE5},
{8'hF7, 8'hF4, 8'hE9},
{8'hFA, 8'hF5, 8'hED},
{8'hF4, 8'hF0, 8'hE8},
{8'hCA, 8'hC6, 8'hBE},
{8'hD3, 8'hD3, 8'hC7},
{8'hEA, 8'hEA, 8'hDE},
{8'hEA, 8'hEB, 8'hDE},
{8'hDA, 8'hDB, 8'hCD},
{8'hA6, 8'hA7, 8'h97},
{8'hCD, 8'hCE, 8'hBD},
{8'hE0, 8'hE1, 8'hD0},
{8'hAF, 8'hB0, 8'h9C},
{8'h93, 8'h94, 8'h70},
{8'hAF, 8'hAF, 8'h8D},
{8'hB7, 8'hB7, 8'h98},
{8'h9E, 8'h9E, 8'h83},
{8'hC9, 8'hC8, 8'hB1},
{8'hEE, 8'hED, 8'hDB},
{8'hF7, 8'hF4, 8'hE5},
{8'hF9, 8'hF7, 8'hEA},
{8'hF2, 8'hF1, 8'hED},
{8'hF2, 8'hF1, 8'hEE},
{8'hF3, 8'hF1, 8'hED},
{8'hEB, 8'hE9, 8'hDE},
{8'hE2, 8'hE0, 8'hC9},
{8'hDD, 8'hDC, 8'hB3},
{8'hD6, 8'hD6, 8'h9C},
{8'hEF, 8'hF1, 8'hB1},
{8'hF0, 8'hF2, 8'hD8},
{8'hEC, 8'hED, 8'hDC},
{8'hEF, 8'hEF, 8'hE3},
{8'hEE, 8'hED, 8'hE8},
{8'hA9, 8'hA8, 8'hA7},
{8'h7C, 8'h7A, 8'h7B},
{8'h7E, 8'h7C, 8'h7D},
{8'h7F, 8'h7E, 8'h7C},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'h80, 8'h7E, 8'h83},
{8'h82, 8'h80, 8'h84},
{8'h79, 8'h77, 8'h7A},
{8'h82, 8'h80, 8'h82},
{8'hB5, 8'hB4, 8'hB4},
{8'hE9, 8'hE8, 8'hE6},
{8'hFA, 8'hF9, 8'hF6},
{8'hF5, 8'hF4, 8'hF0},
{8'hFA, 8'hF9, 8'hFD},
{8'hF9, 8'hF8, 8'hFF},
{8'hF7, 8'hF6, 8'hFC},
{8'hF7, 8'hF7, 8'hF8},
{8'hFB, 8'hFB, 8'hF3},
{8'hF1, 8'hF4, 8'hDE},
{8'hC8, 8'hCE, 8'hAB},
{8'hAC, 8'hB3, 8'h8A},
{8'hDF, 8'hE6, 8'hC9},
{8'hB8, 8'hBC, 8'hA2},
{8'hDF, 8'hDE, 8'hCA},
{8'hF1, 8'hEA, 8'hE0},
{8'hF5, 8'hEB, 8'hDE},
{8'hF3, 8'hEE, 8'hC8},
{8'hE4, 8'hE5, 8'h97},
{8'hD1, 8'hD7, 8'h6E},
{8'hD4, 8'hD9, 8'h97},
{8'hE0, 8'hE4, 8'hB0},
{8'hE3, 8'hE5, 8'hC3},
{8'hE4, 8'hE5, 8'hD3},
{8'hE1, 8'hE3, 8'hD7},
{8'hCE, 8'hD1, 8'hC4},
{8'hD9, 8'hDD, 8'hC9},
{8'hEC, 8'hF2, 8'hD7},
{8'hEB, 8'hF1, 8'hCE},
{8'hE3, 8'hEA, 8'hC6},
{8'hF1, 8'hF7, 8'hDC},
{8'hD5, 8'hD7, 8'hCF},
{8'h13, 8'h12, 8'h20},
{8'h01, 8'h00, 8'h1B},
{8'h07, 8'h04, 8'h22},
{8'h01, 8'h00, 8'h1A},
{8'h0F, 8'h1A, 8'h57},
{8'h21, 8'h4D, 8'h95},
{8'h03, 8'h17, 8'h3C},
{8'h01, 8'h03, 8'h17},
{8'h0D, 8'h3C, 8'h7D},
{8'h0D, 8'h59, 8'hC0},
{8'h10, 8'h54, 8'hBB},
{8'h0D, 8'h52, 8'hB7},
{8'h0D, 8'h58, 8'hAC},
{8'h09, 8'h52, 8'hB5},
{8'h19, 8'h52, 8'hCA},
{8'h29, 8'h46, 8'hA2},
{8'h08, 8'h0D, 8'h2D},
{8'h00, 8'h00, 8'h18},
{8'h0F, 8'h1E, 8'h6B},
{8'h22, 8'h49, 8'hBA},
{8'h16, 8'h48, 8'h9C},
{8'h12, 8'h4F, 8'h9D},
{8'h13, 8'h57, 8'hBE},
{8'h13, 8'h49, 8'hCE},
{8'h28, 8'h4B, 8'hBE},
{8'h17, 8'h2B, 8'h67},
{8'h00, 8'h06, 8'h23},
{8'h00, 8'h05, 8'h29},
{8'h01, 8'h15, 8'h4F},
{8'h26, 8'h3F, 8'h8D},
{8'h1A, 8'h27, 8'h6C},
{8'h00, 8'h00, 8'h24},
{8'h00, 8'h01, 8'h1E},
{8'h01, 8'h00, 8'h28},
{8'h01, 8'h00, 8'h1D},
{8'h00, 8'h00, 8'h00},
{8'h83, 8'h81, 8'h6D},
{8'hF6, 8'hF4, 8'hDC},
{8'hEF, 8'hEC, 8'hD7},
{8'hE5, 8'hE2, 8'hD0},
{8'hD7, 8'hD3, 8'hC6},
{8'hA9, 8'hA5, 8'h9B},
{8'h95, 8'h90, 8'h8B},
{8'h81, 8'h7C, 8'h78},
{8'hCF, 8'hCF, 8'hC4},
{8'hE2, 8'hE2, 8'hD7},
{8'hB7, 8'hB7, 8'hAB},
{8'hE6, 8'hE6, 8'hDB},
{8'hDC, 8'hDC, 8'hCF},
{8'h8E, 8'h8F, 8'h82},
{8'hCF, 8'hD0, 8'hC3},
{8'hFF, 8'hFF, 8'hF2},
{8'hE9, 8'hE9, 8'hD0},
{8'hA3, 8'hA4, 8'h88},
{8'h94, 8'h94, 8'h7A},
{8'hB7, 8'hB6, 8'h9F},
{8'hED, 8'hEC, 8'hDA},
{8'hFC, 8'hFA, 8'hEE},
{8'hF3, 8'hF0, 8'hEA},
{8'hC8, 8'hC5, 8'hC3},
{8'hD9, 8'hD6, 8'hDC},
{8'hF0, 8'hEE, 8'hF2},
{8'hF1, 8'hEF, 8'hED},
{8'hF4, 8'hF2, 8'hE2},
{8'hE6, 8'hE6, 8'hC3},
{8'hD7, 8'hD9, 8'h9D},
{8'hD1, 8'hD6, 8'h83},
{8'hCF, 8'hD5, 8'h7B},
{8'hE6, 8'hE8, 8'hCF},
{8'hEC, 8'hED, 8'hDF},
{8'hF3, 8'hF3, 8'hEA},
{8'hF4, 8'hF3, 8'hF0},
{8'hF6, 8'hF4, 8'hF5},
{8'hDD, 8'hDB, 8'hDC},
{8'h9E, 8'h9C, 8'h9C},
{8'h7B, 8'h7A, 8'h77},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'h7C, 8'h7A, 8'h7F},
{8'h7C, 8'h7A, 8'h7E},
{8'h80, 8'h7E, 8'h81},
{8'h7B, 8'h79, 8'h7B},
{8'h78, 8'h76, 8'h76},
{8'hA3, 8'hA2, 8'hA0},
{8'hD4, 8'hD3, 8'hD0},
{8'hF1, 8'hF0, 8'hEB},
{8'hF8, 8'hF9, 8'hEE},
{8'hFB, 8'hFC, 8'hF5},
{8'hFF, 8'hFF, 8'hFD},
{8'hFB, 8'hFB, 8'hFB},
{8'hF3, 8'hF4, 8'hEF},
{8'hE2, 8'hE4, 8'hD5},
{8'hAB, 8'hAF, 8'h94},
{8'hA2, 8'hA9, 8'h86},
{8'h95, 8'hA1, 8'h90},
{8'h97, 8'hA0, 8'h8D},
{8'hE9, 8'hEA, 8'hD9},
{8'hF3, 8'hEF, 8'hE3},
{8'hF8, 8'hF0, 8'hE8},
{8'hFB, 8'hF6, 8'hE1},
{8'hF5, 8'hF6, 8'hC7},
{8'hEB, 8'hF2, 8'hAF},
{8'hE7, 8'hEB, 8'hBA},
{8'hE3, 8'hE6, 8'hC0},
{8'hF1, 8'hF3, 8'hDB},
{8'hF3, 8'hF4, 8'hE7},
{8'hEE, 8'hF1, 8'hE6},
{8'hE4, 8'hE8, 8'hD8},
{8'hE8, 8'hEE, 8'hD4},
{8'hE9, 8'hF3, 8'hD1},
{8'hDF, 8'hE9, 8'hBB},
{8'hE4, 8'hEE, 8'hBE},
{8'hEF, 8'hF6, 8'hD2},
{8'h82, 8'h85, 8'h7D},
{8'h02, 8'h01, 8'h17},
{8'h05, 8'h03, 8'h26},
{8'h03, 8'h01, 8'h1C},
{8'h03, 8'h01, 8'h15},
{8'h15, 8'h2C, 8'h74},
{8'h1B, 8'h54, 8'hA7},
{8'h08, 8'h1F, 8'h51},
{8'h02, 8'h04, 8'h25},
{8'h18, 8'h40, 8'h8B},
{8'h0F, 8'h54, 8'hC0},
{8'h14, 8'h54, 8'hBA},
{8'h11, 8'h52, 8'hB3},
{8'h16, 8'h52, 8'hAF},
{8'h13, 8'h54, 8'hA8},
{8'h1C, 8'h53, 8'hB9},
{8'h22, 8'h40, 8'h99},
{8'h03, 8'h09, 8'h2E},
{8'h05, 8'h0A, 8'h37},
{8'h1E, 8'h3A, 8'h9B},
{8'h1B, 8'h51, 8'hBD},
{8'h12, 8'h4E, 8'hA2},
{8'h13, 8'h4A, 8'hA2},
{8'h1C, 8'h50, 8'hB7},
{8'h14, 8'h4E, 8'hC5},
{8'h10, 8'h4F, 8'hC6},
{8'h19, 8'h4D, 8'hAA},
{8'h06, 8'h1B, 8'h4D},
{8'h02, 8'h05, 8'h18},
{8'h01, 8'h06, 8'h25},
{8'h06, 8'h09, 8'h42},
{8'h11, 8'h15, 8'h50},
{8'h03, 8'h04, 8'h23},
{8'h00, 8'h01, 8'h16},
{8'h01, 8'h00, 8'h25},
{8'h00, 8'h01, 8'h25},
{8'h00, 8'h00, 8'h0B},
{8'h33, 8'h2F, 8'h2D},
{8'hEC, 8'hE7, 8'hDF},
{8'hF5, 8'hF1, 8'hE4},
{8'hF0, 8'hEC, 8'hDD},
{8'hE3, 8'hE0, 8'hD2},
{8'h99, 8'h95, 8'h8B},
{8'h7B, 8'h76, 8'h72},
{8'h81, 8'h7C, 8'h7B},
{8'hDE, 8'hDE, 8'hD6},
{8'hCF, 8'hD0, 8'hC6},
{8'h74, 8'h74, 8'h6B},
{8'hD6, 8'hD5, 8'hCE},
{8'hFF, 8'hFF, 8'hFB},
{8'hCE, 8'hCE, 8'hC7},
{8'h7D, 8'h7D, 8'h76},
{8'hD7, 8'hD7, 8'hD1},
{8'hFF, 8'hFF, 8'hF5},
{8'hF4, 8'hF4, 8'hE6},
{8'hC7, 8'hC8, 8'hB7},
{8'hD0, 8'hD1, 8'hC1},
{8'hF6, 8'hF6, 8'hE9},
{8'hE6, 8'hE5, 8'hDE},
{8'hA0, 8'h9F, 8'h9E},
{8'h77, 8'h75, 8'h78},
{8'h87, 8'h85, 8'h87},
{8'hB5, 8'hB3, 8'hB4},
{8'hEE, 8'hEC, 8'hE9},
{8'hF1, 8'hEF, 8'hE3},
{8'hF5, 8'hF4, 8'hD8},
{8'hE7, 8'hE8, 8'hB7},
{8'hCF, 8'hD1, 8'h8E},
{8'hDA, 8'hDE, 8'h93},
{8'hEE, 8'hF0, 8'hDC},
{8'hF6, 8'hF7, 8'hEB},
{8'hFB, 8'hFB, 8'hF5},
{8'hF7, 8'hF6, 8'hF4},
{8'hF2, 8'hF0, 8'hF1},
{8'hF4, 8'hF2, 8'hF3},
{8'hE6, 8'hE4, 8'hE3},
{8'h82, 8'h81, 8'h7D},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'h83, 8'h81, 8'h86},
{8'h80, 8'h7E, 8'h82},
{8'h7B, 8'h79, 8'h7C},
{8'h83, 8'h81, 8'h83},
{8'h82, 8'h81, 8'h80},
{8'h7A, 8'h79, 8'h78},
{8'h84, 8'h82, 8'h80},
{8'hDD, 8'hDC, 8'hD5},
{8'hEA, 8'hF1, 8'hC2},
{8'hEA, 8'hF1, 8'hC9},
{8'hFC, 8'hFE, 8'hEB},
{8'hF4, 8'hF5, 8'hF0},
{8'hF3, 8'hF2, 8'hF5},
{8'h98, 8'h98, 8'h99},
{8'h7E, 8'h80, 8'h78},
{8'h8A, 8'h8E, 8'h81},
{8'h83, 8'h92, 8'h8F},
{8'hCC, 8'hD9, 8'hCE},
{8'hF8, 8'hFD, 8'hED},
{8'hFC, 8'hFC, 8'hEF},
{8'hFE, 8'hFB, 8'hF8},
{8'hFB, 8'hF7, 8'hF4},
{8'hF0, 8'hF1, 8'hE1},
{8'hE8, 8'hEE, 8'hD1},
{8'hE9, 8'hED, 8'hCE},
{8'hF2, 8'hF3, 8'hDC},
{8'hFA, 8'hFB, 8'hEE},
{8'hF8, 8'hF9, 8'hF3},
{8'hF5, 8'hF7, 8'hF0},
{8'hE3, 8'hE8, 8'hD7},
{8'hE1, 8'hEB, 8'hCA},
{8'hE3, 8'hEF, 8'hC3},
{8'hE1, 8'hED, 8'hB8},
{8'hE8, 8'hF4, 8'hBB},
{8'hDC, 8'hE6, 8'hBA},
{8'h22, 8'h27, 8'h20},
{8'h01, 8'h01, 8'h1A},
{8'h01, 8'h00, 8'h2A},
{8'h04, 8'h04, 8'h1E},
{8'h02, 8'h04, 8'h10},
{8'h18, 8'h3E, 8'h92},
{8'h15, 8'h55, 8'hBA},
{8'h0C, 8'h29, 8'h70},
{8'h04, 8'h04, 8'h38},
{8'h23, 8'h42, 8'hA1},
{8'h12, 8'h4E, 8'hC7},
{8'h1B, 8'h52, 8'hBC},
{8'h16, 8'h4F, 8'hB2},
{8'h1C, 8'h4B, 8'hC1},
{8'h17, 8'h55, 8'hAC},
{8'h18, 8'h56, 8'hB7},
{8'h15, 8'h3E, 8'h9A},
{8'h00, 8'h09, 8'h39},
{8'h11, 8'h23, 8'h63},
{8'h1F, 8'h4C, 8'hB3},
{8'h0E, 8'h58, 8'hB4},
{8'h0C, 8'h51, 8'hB5},
{8'h15, 8'h42, 8'hAE},
{8'h24, 8'h4A, 8'hAA},
{8'h17, 8'h56, 8'hA9},
{8'h01, 8'h5A, 8'hBF},
{8'h08, 8'h57, 8'hCD},
{8'h17, 8'h3A, 8'h8C},
{8'h0B, 8'h06, 8'h1A},
{8'h05, 8'h03, 8'h0C},
{8'h05, 8'h00, 8'h2A},
{8'h07, 8'h02, 8'h33},
{8'h06, 8'h03, 8'h1A},
{8'h01, 8'h02, 8'h10},
{8'h00, 8'h01, 8'h22},
{8'h00, 8'h00, 8'h29},
{8'h01, 8'h03, 8'h1B},
{8'h02, 8'h01, 8'h05},
{8'h9E, 8'h99, 8'h9C},
{8'hFC, 8'hFA, 8'hF6},
{8'hF5, 8'hF0, 8'hE4},
{8'hF8, 8'hF5, 8'hE7},
{8'hC1, 8'hBD, 8'hB2},
{8'h7C, 8'h77, 8'h73},
{8'h84, 8'h7E, 8'h7F},
{8'hE0, 8'hDF, 8'hDA},
{8'hE5, 8'hE4, 8'hDF},
{8'h7D, 8'h7D, 8'h78},
{8'h9B, 8'h9A, 8'h96},
{8'hF9, 8'hF8, 8'hF5},
{8'hFF, 8'hFE, 8'hFC},
{8'hAF, 8'hAE, 8'hAD},
{8'h84, 8'h82, 8'h82},
{8'hDF, 8'hDD, 8'hDD},
{8'hFD, 8'hFC, 8'hF9},
{8'hFD, 8'hFD, 8'hF5},
{8'hB8, 8'hB8, 8'hAD},
{8'h88, 8'h88, 8'h7E},
{8'h82, 8'h81, 8'h7D},
{8'h78, 8'h76, 8'h79},
{8'h83, 8'h80, 8'h87},
{8'h7E, 8'h7E, 8'h72},
{8'h81, 8'h81, 8'h76},
{8'hDA, 8'hD8, 8'hD3},
{8'hEF, 8'hEB, 8'hE7},
{8'hDB, 8'hD7, 8'hCF},
{8'hED, 8'hEA, 8'hD8},
{8'hE6, 8'hE2, 8'hC5},
{8'hED, 8'hEB, 8'hC8},
{8'hF3, 8'hF3, 8'hE3},
{8'hF1, 8'hF1, 8'hE6},
{8'hD2, 8'hD1, 8'hCC},
{8'hA6, 8'hA5, 8'hA5},
{8'hA1, 8'h9F, 8'hA2},
{8'hA6, 8'hA4, 8'hA5},
{8'h9C, 8'h9A, 8'h98},
{8'h7D, 8'h7C, 8'h77},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'h7F, 8'h7C, 8'h82},
{8'h7E, 8'h7C, 8'h81},
{8'hFF, 8'hD7, 8'h00},
{8'h7F, 8'h7D, 8'h7E},
{8'h7E, 8'h7D, 8'h7A},
{8'h80, 8'h7F, 8'h7A},
{8'h7A, 8'h79, 8'h72},
{8'hAE, 8'hAE, 8'hA4},
{8'hD1, 8'hD7, 8'hB4},
{8'hE6, 8'hEB, 8'hCB},
{8'hE9, 8'hED, 8'hD8},
{8'hDE, 8'hE0, 8'hD5},
{8'hC0, 8'hC1, 8'hBE},
{8'h7C, 8'h7B, 8'h7D},
{8'h7C, 8'h7C, 8'h7E},
{8'h7C, 8'h7C, 8'h7E},
{8'h81, 8'h89, 8'h8E},
{8'hF1, 8'hF5, 8'hF5},
{8'hFC, 8'hFD, 8'hF7},
{8'hFB, 8'hFA, 8'hF5},
{8'hF9, 8'hF7, 8'hF4},
{8'hF0, 8'hEE, 8'hEC},
{8'hED, 8'hEE, 8'hE7},
{8'hE8, 8'hEB, 8'hDD},
{8'hEC, 8'hF2, 8'hD1},
{8'hEA, 8'hEE, 8'hD2},
{8'hE9, 8'hEE, 8'hD7},
{8'hF2, 8'hF7, 8'hE1},
{8'hEF, 8'hF7, 8'hD7},
{8'hE3, 8'hEE, 8'hC6},
{8'hE0, 8'hED, 8'hC2},
{8'hE2, 8'hF0, 8'hC4},
{8'hDE, 8'hF3, 8'hB9},
{8'hE4, 8'hFA, 8'hCB},
{8'h8F, 8'h9E, 8'h85},
{8'h00, 8'h02, 8'h02},
{8'h04, 8'h03, 8'h19},
{8'h03, 8'h03, 8'h22},
{8'h01, 8'h03, 8'h1C},
{8'h0C, 8'h10, 8'h25},
{8'h16, 8'h4C, 8'hAC},
{8'h15, 8'h56, 8'hC0},
{8'h11, 8'h38, 8'h8E},
{8'h03, 8'h09, 8'h53},
{8'h22, 8'h44, 8'hA2},
{8'h1A, 8'h4E, 8'hBB},
{8'h1A, 8'h52, 8'hBB},
{8'h12, 8'h50, 8'hB8},
{8'h18, 8'h4F, 8'hC6},
{8'h18, 8'h56, 8'hB4},
{8'h19, 8'h54, 8'hB0},
{8'h0C, 8'h39, 8'h91},
{8'h01, 8'h13, 8'h57},
{8'h16, 8'h40, 8'h91},
{8'h19, 8'h52, 8'hB9},
{8'h0D, 8'h57, 8'hB7},
{8'h0F, 8'h50, 8'hB8},
{8'h12, 8'h43, 8'hAF},
{8'h1F, 8'h4C, 8'hAB},
{8'h16, 8'h56, 8'hA7},
{8'h0B, 8'h5A, 8'hB9},
{8'h0A, 8'h57, 8'hC9},
{8'h1D, 8'h52, 8'hB5},
{8'h0D, 8'h24, 8'h62},
{8'h05, 8'h03, 8'h1B},
{8'h05, 8'h01, 8'h1E},
{8'h0B, 8'h01, 8'h1F},
{8'h0D, 8'h06, 8'h17},
{8'h04, 8'h03, 8'h15},
{8'h00, 8'h01, 8'h22},
{8'h00, 8'h01, 8'h27},
{8'h02, 8'h03, 8'h22},
{8'h01, 8'h01, 8'h11},
{8'h34, 8'h30, 8'h3E},
{8'hEF, 8'hED, 8'hF2},
{8'hFA, 8'hF7, 8'hF2},
{8'hFD, 8'hFC, 8'hF5},
{8'hE4, 8'hE2, 8'hDB},
{8'h7E, 8'h7B, 8'h77},
{8'h7F, 8'h7B, 8'h7B},
{8'hE8, 8'hE6, 8'hE2},
{8'hF0, 8'hEE, 8'hEB},
{8'h85, 8'h84, 8'h82},
{8'h7C, 8'h7A, 8'h7A},
{8'hD5, 8'hD3, 8'hD5},
{8'hFF, 8'hFF, 8'hFF},
{8'hEA, 8'hE9, 8'hE8},
{8'h82, 8'h81, 8'h80},
{8'h8C, 8'h8A, 8'h8E},
{8'hE1, 8'hDF, 8'hDF},
{8'hFE, 8'hFE, 8'hF8},
{8'hF8, 8'hF8, 8'hEF},
{8'hA1, 8'hA1, 8'h97},
{8'h7A, 8'h79, 8'h75},
{8'h83, 8'h81, 8'h83},
{8'h7A, 8'h77, 8'h7D},
{8'h91, 8'h91, 8'h89},
{8'hD2, 8'hD2, 8'hCC},
{8'hEC, 8'hEA, 8'hE8},
{8'hAE, 8'hAB, 8'hAC},
{8'h89, 8'h86, 8'h87},
{8'hE7, 8'hE3, 8'hE1},
{8'hF9, 8'hF5, 8'hF0},
{8'hFB, 8'hF8, 8'hF0},
{8'hF9, 8'hF8, 8'hF0},
{8'hF9, 8'hF8, 8'hF2},
{8'hD7, 8'hD6, 8'hD3},
{8'h7A, 8'h78, 8'h78},
{8'h7C, 8'h7A, 8'h7C},
{8'h7B, 8'h79, 8'h7B},
{8'h7B, 8'h79, 8'h7A},
{8'h80, 8'h7F, 8'h7F},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'h7F, 8'h7C, 8'h83},
{8'h7F, 8'h7C, 8'h82},
{8'hFF, 8'hD7, 8'h00},
{8'h7F, 8'h7E, 8'h7D},
{8'h7F, 8'h7F, 8'h79},
{8'h7E, 8'h7E, 8'h75},
{8'h8E, 8'h8E, 8'h82},
{8'h95, 8'h95, 8'h89},
{8'h7B, 8'h7C, 8'h78},
{8'hD6, 8'hD7, 8'hD2},
{8'hE2, 8'hE4, 8'hDA},
{8'hCF, 8'hD2, 8'hC5},
{8'h8A, 8'h8C, 8'h81},
{8'h7F, 8'h80, 8'h7A},
{8'h7A, 8'h7A, 8'h79},
{8'h7C, 8'h7C, 8'h7F},
{8'h7E, 8'h7A, 8'h81},
{8'hEE, 8'hEC, 8'hF0},
{8'hFE, 8'hFD, 8'hFF},
{8'hF9, 8'hF7, 8'hF8},
{8'hF3, 8'hF3, 8'hEE},
{8'hF3, 8'hF3, 8'hEA},
{8'hE4, 8'hE4, 8'hD9},
{8'hCF, 8'hCF, 8'hC1},
{8'hC7, 8'hCF, 8'hA8},
{8'hD4, 8'hDB, 8'hB9},
{8'hE6, 8'hEF, 8'hCE},
{8'hE1, 8'hED, 8'hC1},
{8'hE1, 8'hF0, 8'hB5},
{8'hE1, 8'hF2, 8'hB3},
{8'hE0, 8'hF1, 8'hBD},
{8'hDF, 8'hEE, 8'hC5},
{8'hE3, 8'hF6, 8'hC0},
{8'hDD, 8'hF0, 8'hD5},
{8'h3F, 8'h48, 8'h4C},
{8'h00, 8'h00, 8'h0A},
{8'h04, 8'h01, 8'h15},
{8'h00, 8'h02, 8'h1A},
{8'h00, 8'h03, 8'h23},
{8'h13, 8'h19, 8'h44},
{8'h13, 8'h55, 8'hBB},
{8'h16, 8'h55, 8'hB9},
{8'h16, 8'h47, 8'hA2},
{8'h03, 8'h18, 8'h6D},
{8'h1C, 8'h45, 8'h98},
{8'h1F, 8'h51, 8'hAA},
{8'h16, 8'h54, 8'hB8},
{8'h0C, 8'h53, 8'hBD},
{8'h11, 8'h55, 8'hBD},
{8'h19, 8'h56, 8'hB6},
{8'h19, 8'h4E, 8'hA5},
{8'h11, 8'h32, 8'h83},
{8'h05, 8'h29, 8'h7E},
{8'h18, 8'h4E, 8'hAB},
{8'h16, 8'h52, 8'hB9},
{8'h14, 8'h54, 8'hC3},
{8'h16, 8'h50, 8'hB1},
{8'h0E, 8'h48, 8'hA9},
{8'h14, 8'h51, 8'hB4},
{8'h14, 8'h51, 8'hB4},
{8'h16, 8'h52, 8'hB7},
{8'h12, 8'h51, 8'hB4},
{8'h16, 8'h58, 8'hBE},
{8'h07, 8'h44, 8'hAB},
{8'h04, 8'h0D, 8'h42},
{8'h02, 8'h00, 8'h20},
{8'h0B, 8'h01, 8'h16},
{8'h0B, 8'h02, 8'h13},
{8'h03, 8'h02, 8'h1B},
{8'h00, 8'h03, 8'h23},
{8'h00, 8'h02, 8'h24},
{8'h04, 8'h00, 8'h21},
{8'h00, 8'h00, 8'h19},
{8'h03, 8'h03, 8'h14},
{8'hAA, 8'hAA, 8'hB4},
{8'hFB, 8'hFC, 8'hFE},
{8'hFC, 8'hFB, 8'hFB},
{8'hE9, 8'hE8, 8'hE5},
{8'h81, 8'h7F, 8'h7C},
{8'h86, 8'h82, 8'h81},
{8'hEF, 8'hEE, 8'hE8},
{8'hFA, 8'hF9, 8'hF5},
{8'h8D, 8'h8C, 8'h8C},
{8'h77, 8'h75, 8'h78},
{8'h97, 8'h95, 8'h98},
{8'hF4, 8'hF3, 8'hF2},
{8'hFD, 8'hFC, 8'hF7},
{8'hAE, 8'hAE, 8'hA8},
{8'h72, 8'h70, 8'h73},
{8'h88, 8'h86, 8'h86},
{8'hD5, 8'hD5, 8'hCF},
{8'hFF, 8'hFF, 8'hF6},
{8'hEC, 8'hEC, 8'hE2},
{8'h91, 8'h90, 8'h8A},
{8'h77, 8'h76, 8'h75},
{8'h80, 8'h7E, 8'h82},
{8'h7D, 8'h7B, 8'h81},
{8'hB2, 8'hAF, 8'hB4},
{8'hAE, 8'hAC, 8'hAF},
{8'h74, 8'h72, 8'h74},
{8'hA5, 8'hA4, 8'hA3},
{8'hFB, 8'hFB, 8'hF9},
{8'hF3, 8'hF2, 8'hEF},
{8'hFA, 8'hFA, 8'hF6},
{8'hE8, 8'hE7, 8'hE4},
{8'hF6, 8'hF5, 8'hF2},
{8'hF0, 8'hEF, 8'hED},
{8'h93, 8'h92, 8'h91},
{8'h7C, 8'h7A, 8'h7C},
{8'hFF, 8'hD7, 8'h00},
{8'h7F, 8'h7D, 8'h81},
{8'h7F, 8'h7D, 8'h82},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'h7F, 8'h7C, 8'h83},
{8'h7F, 8'h7D, 8'h82},
{8'hFF, 8'hD7, 8'h00},
{8'h7F, 8'h7D, 8'h7D},
{8'h7D, 8'h7D, 8'h78},
{8'h88, 8'h87, 8'h81},
{8'h94, 8'h94, 8'h8B},
{8'h7A, 8'h7A, 8'h70},
{8'h92, 8'h93, 8'h8E},
{8'hDB, 8'hDC, 8'hD6},
{8'hE6, 8'hE7, 8'hDE},
{8'hD7, 8'hD9, 8'hCE},
{8'hAE, 8'hB0, 8'hA6},
{8'h80, 8'h81, 8'h7B},
{8'h7B, 8'h7B, 8'h7A},
{8'h7D, 8'h7C, 8'h80},
{8'h7D, 8'h7A, 8'h81},
{8'hBA, 8'hB8, 8'hBD},
{8'hF9, 8'hF8, 8'hF9},
{8'hFC, 8'hFC, 8'hFB},
{8'hF9, 8'hF8, 8'hF4},
{8'hDF, 8'hDE, 8'hD8},
{8'h9A, 8'h9A, 8'h91},
{8'h7C, 8'h7C, 8'h70},
{8'h7B, 8'h80, 8'h67},
{8'h7F, 8'h84, 8'h70},
{8'hA2, 8'hA9, 8'h93},
{8'hD5, 8'hE0, 8'hBC},
{8'hE4, 8'hF2, 8'hBE},
{8'hE1, 8'hF2, 8'hB6},
{8'hE0, 8'hF1, 8'hBC},
{8'hE3, 8'hF1, 8'hC5},
{8'hED, 8'hE9, 8'hBC},
{8'h78, 8'h6E, 8'h58},
{8'h12, 8'h06, 8'h0D},
{8'h0B, 8'h03, 8'h1A},
{8'h06, 8'h01, 8'h21},
{8'h00, 8'h01, 8'h25},
{8'h00, 8'h00, 8'h2F},
{8'h16, 8'h26, 8'h63},
{8'h14, 8'h55, 8'hBC},
{8'h12, 8'h51, 8'hB5},
{8'h1B, 8'h50, 8'hAC},
{8'h0A, 8'h28, 8'h7D},
{8'h1B, 8'h43, 8'h98},
{8'h1D, 8'h52, 8'hAD},
{8'h16, 8'h54, 8'hB8},
{8'h0D, 8'h53, 8'hBC},
{8'h10, 8'h52, 8'hBA},
{8'h15, 8'h52, 8'hB3},
{8'h1B, 8'h50, 8'hA9},
{8'h09, 8'h2E, 8'h81},
{8'h17, 8'h46, 8'h9A},
{8'h1C, 8'h52, 8'hAF},
{8'h14, 8'h50, 8'hB7},
{8'h15, 8'h55, 8'hC3},
{8'h16, 8'h50, 8'hB2},
{8'h0E, 8'h48, 8'hA9},
{8'h15, 8'h51, 8'hB3},
{8'h14, 8'h51, 8'hB3},
{8'h17, 8'h55, 8'hB9},
{8'h11, 8'h51, 8'hB5},
{8'h17, 8'h56, 8'hBD},
{8'h19, 8'h57, 8'hBB},
{8'h15, 8'h2F, 8'h6F},
{8'h00, 8'h02, 8'h31},
{8'h05, 8'h04, 8'h22},
{8'h04, 8'h01, 8'h17},
{8'h02, 8'h02, 8'h1C},
{8'h00, 8'h03, 8'h22},
{8'h01, 8'h01, 8'h23},
{8'h05, 8'h00, 8'h20},
{8'h01, 8'h01, 8'h1A},
{8'h01, 8'h00, 8'h14},
{8'h44, 8'h43, 8'h50},
{8'hFE, 8'hFD, 8'hFE},
{8'hFF, 8'hFF, 8'hFF},
{8'hC8, 8'hC8, 8'hC5},
{8'h79, 8'h77, 8'h75},
{8'h98, 8'h95, 8'h93},
{8'hF6, 8'hF6, 8'hF0},
{8'hFB, 8'hFB, 8'hF6},
{8'h96, 8'h95, 8'h94},
{8'hFF, 8'hD7, 8'h00},
{8'h7C, 8'h7A, 8'h7D},
{8'hBC, 8'hBB, 8'hBB},
{8'hFE, 8'hFD, 8'hF9},
{8'hDB, 8'hDB, 8'hD5},
{8'h81, 8'h7F, 8'h81},
{8'h79, 8'h78, 8'h77},
{8'h83, 8'h82, 8'h7D},
{8'hB7, 8'hB6, 8'hAF},
{8'hF4, 8'hF4, 8'hED},
{8'hDA, 8'hD9, 8'hD4},
{8'h7D, 8'h7B, 8'h7B},
{8'h7D, 8'h7B, 8'h7E},
{8'h7E, 8'h7C, 8'h81},
{8'h7E, 8'h7C, 8'h80},
{8'h7D, 8'h7B, 8'h7E},
{8'h7B, 8'h79, 8'h7B},
{8'hCC, 8'hCB, 8'hCA},
{8'hFD, 8'hFD, 8'hFB},
{8'hF6, 8'hF5, 8'hF2},
{8'hEF, 8'hEF, 8'hEB},
{8'h95, 8'h94, 8'h90},
{8'hD8, 8'hD7, 8'hD4},
{8'hF6, 8'hF5, 8'hF3},
{8'hB3, 8'hB1, 8'hB1},
{8'h79, 8'h77, 8'h79},
{8'hFF, 8'hD7, 8'h00},
{8'h7F, 8'h7D, 8'h81},
{8'h7F, 8'h7D, 8'h82},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'h7F, 8'h7D, 8'h82},
{8'h7F, 8'h7D, 8'h82},
{8'hFF, 8'hD7, 8'h00},
{8'h7E, 8'h7C, 8'h7D},
{8'h7C, 8'h7B, 8'h78},
{8'h8F, 8'h8E, 8'h89},
{8'h84, 8'h83, 8'h7E},
{8'h7D, 8'h7D, 8'h76},
{8'h87, 8'h88, 8'h85},
{8'hDE, 8'hDF, 8'hDA},
{8'hF9, 8'hF9, 8'hF4},
{8'hED, 8'hEE, 8'hE5},
{8'hB7, 8'hB8, 8'hB0},
{8'h7F, 8'h7F, 8'h7B},
{8'h81, 8'h81, 8'h82},
{8'h80, 8'h7F, 8'h83},
{8'h7F, 8'h7D, 8'h82},
{8'h7F, 8'h7D, 8'h82},
{8'h98, 8'h96, 8'h99},
{8'hCA, 8'hC9, 8'hC9},
{8'hBE, 8'hBD, 8'hBA},
{8'h87, 8'h86, 8'h82},
{8'h7B, 8'h7B, 8'h75},
{8'h82, 8'h81, 8'h7B},
{8'h7E, 8'h80, 8'h78},
{8'h7C, 8'h7E, 8'h79},
{8'h79, 8'h7D, 8'h74},
{8'hC6, 8'hCE, 8'hB4},
{8'hE6, 8'hF3, 8'hC3},
{8'hE1, 8'hF2, 8'hB6},
{8'hE0, 8'hF2, 8'hBA},
{8'hE6, 8'hF3, 8'hC4},
{8'hB6, 8'h96, 8'h6A},
{8'h72, 8'h44, 8'h28},
{8'h37, 8'h11, 8'h10},
{8'h10, 8'h00, 8'h16},
{8'h08, 8'h01, 8'h25},
{8'h02, 8'h02, 8'h26},
{8'h00, 8'h01, 8'h34},
{8'h1B, 8'h39, 8'h83},
{8'h11, 8'h52, 8'hBA},
{8'h16, 8'h54, 8'hB9},
{8'h1C, 8'h52, 8'hB0},
{8'h11, 8'h3A, 8'h92},
{8'h17, 8'h46, 8'h9D},
{8'h1C, 8'h51, 8'hAF},
{8'h16, 8'h54, 8'hB8},
{8'h0E, 8'h52, 8'hBB},
{8'h11, 8'h52, 8'hB9},
{8'h16, 8'h53, 8'hB5},
{8'h18, 8'h4E, 8'hA9},
{8'h0E, 8'h3C, 8'h93},
{8'h1F, 8'h53, 8'hAB},
{8'h1B, 8'h52, 8'hB1},
{8'h16, 8'h52, 8'hBA},
{8'h12, 8'h51, 8'hBE},
{8'h16, 8'h50, 8'hB2},
{8'h0E, 8'h48, 8'hA9},
{8'h15, 8'h51, 8'hB3},
{8'h13, 8'h50, 8'hB3},
{8'h14, 8'h53, 8'hB7},
{8'h14, 8'h54, 8'hB8},
{8'h13, 8'h53, 8'hB9},
{8'h14, 8'h53, 8'hB9},
{8'h1F, 8'h4E, 8'hA0},
{8'h09, 8'h21, 8'h60},
{8'h00, 8'h03, 8'h2D},
{8'h03, 8'h04, 8'h21},
{8'h01, 8'h02, 8'h20},
{8'h00, 8'h03, 8'h21},
{8'h02, 8'h01, 8'h20},
{8'h06, 8'h00, 8'h1D},
{8'h04, 8'h04, 8'h1E},
{8'h04, 8'h04, 8'h18},
{8'h08, 8'h08, 8'h16},
{8'h9F, 8'h9E, 8'hA5},
{8'hCD, 8'hCC, 8'hCD},
{8'h8C, 8'h8A, 8'h8A},
{8'h7A, 8'h77, 8'h77},
{8'hA1, 8'h9D, 8'h9D},
{8'hFA, 8'hFA, 8'hF4},
{8'hF9, 8'hF8, 8'hF3},
{8'h99, 8'h98, 8'h97},
{8'h7D, 8'h7B, 8'h7E},
{8'h7C, 8'h7A, 8'h7D},
{8'h83, 8'h81, 8'h81},
{8'hCD, 8'hCC, 8'hC8},
{8'hF5, 8'hF5, 8'hEF},
{8'h95, 8'h93, 8'h95},
{8'h81, 8'h7F, 8'h80},
{8'h7F, 8'h7D, 8'h7C},
{8'h7B, 8'h7A, 8'h76},
{8'h94, 8'h93, 8'h8F},
{8'hAF, 8'hAE, 8'hAC},
{8'h85, 8'h83, 8'h84},
{8'h83, 8'h81, 8'h84},
{8'h7D, 8'h7B, 8'h80},
{8'h80, 8'h7E, 8'h82},
{8'h7E, 8'h7C, 8'h7F},
{8'h82, 8'h80, 8'h82},
{8'hE1, 8'hE0, 8'hDF},
{8'hF5, 8'hF4, 8'hF2},
{8'hFB, 8'hFA, 8'hF7},
{8'hBC, 8'hBB, 8'hB7},
{8'h7A, 8'h79, 8'h74},
{8'h8F, 8'h8E, 8'h8B},
{8'hEC, 8'hEC, 8'hEA},
{8'hCD, 8'hCC, 8'hCB},
{8'h7D, 8'h7B, 8'h7D},
{8'h7E, 8'h7C, 8'h7F},
{8'h7F, 8'h7D, 8'h81},
{8'h7F, 8'h7D, 8'h82},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'h7F, 8'h7D, 8'h82},
{8'h7F, 8'h7D, 8'h81},
{8'hFF, 8'hD7, 8'h00},
{8'h7F, 8'h7D, 8'h7E},
{8'h80, 8'h7E, 8'h7E},
{8'h7F, 8'h7E, 8'h7C},
{8'h83, 8'h82, 8'h7F},
{8'h81, 8'h80, 8'h7D},
{8'h76, 8'h76, 8'h75},
{8'hB5, 8'hB6, 8'hB1},
{8'hF6, 8'hF7, 8'hF1},
{8'hAC, 8'hAD, 8'hA5},
{8'h73, 8'h75, 8'h6E},
{8'h7E, 8'h7F, 8'h7B},
{8'h7F, 8'h7F, 8'h81},
{8'h7F, 8'h7E, 8'h83},
{8'h82, 8'h80, 8'h85},
{8'h80, 8'h7E, 8'h81},
{8'h7A, 8'h78, 8'h7B},
{8'h80, 8'h7E, 8'h80},
{8'h7A, 8'h78, 8'h78},
{8'h7C, 8'h7B, 8'h79},
{8'h7C, 8'h7B, 8'h78},
{8'h7D, 8'h7C, 8'h79},
{8'h7E, 8'h7F, 8'h81},
{8'h7C, 8'h7D, 8'h82},
{8'h79, 8'h7C, 8'h7C},
{8'hB3, 8'hBB, 8'hA6},
{8'hE6, 8'hF3, 8'hC4},
{8'hE1, 8'hF2, 8'hB6},
{8'hE1, 8'hF4, 8'hBA},
{8'hE2, 8'hEE, 8'hBC},
{8'hAC, 8'h78, 8'h44},
{8'hA4, 8'h5A, 8'h2C},
{8'h84, 8'h45, 8'h33},
{8'h22, 8'h09, 8'h19},
{8'h06, 8'h01, 8'h1E},
{8'h04, 8'h02, 8'h1B},
{8'h02, 8'h04, 8'h31},
{8'h19, 8'h43, 8'h90},
{8'h10, 8'h53, 8'hBA},
{8'h17, 8'h55, 8'hBA},
{8'h19, 8'h50, 8'hAF},
{8'h14, 8'h47, 8'hA1},
{8'h16, 8'h48, 8'hA3},
{8'h1A, 8'h51, 8'hB1},
{8'h14, 8'h52, 8'hB7},
{8'h10, 8'h52, 8'hBA},
{8'h13, 8'h52, 8'hB9},
{8'h17, 8'h54, 8'hB5},
{8'h0F, 8'h49, 8'hA6},
{8'h17, 8'h4F, 8'hA8},
{8'h1A, 8'h51, 8'hAC},
{8'h18, 8'h52, 8'hB2},
{8'h16, 8'h52, 8'hBB},
{8'h11, 8'h4F, 8'hBB},
{8'h16, 8'h50, 8'hB2},
{8'h10, 8'h4A, 8'hAC},
{8'h14, 8'h50, 8'hB2},
{8'h14, 8'h51, 8'hB3},
{8'h13, 8'h51, 8'hB5},
{8'h15, 8'h55, 8'hB9},
{8'h12, 8'h51, 8'hB7},
{8'h0F, 8'h4F, 8'hB6},
{8'h18, 8'h54, 8'hB5},
{8'h1D, 8'h46, 8'h93},
{8'h08, 8'h10, 8'h44},
{8'h02, 8'h03, 8'h26},
{8'h00, 8'h01, 8'h20},
{8'h00, 8'h02, 8'h21},
{8'h04, 8'h01, 8'h1F},
{8'h06, 8'h00, 8'h1A},
{8'h04, 8'h03, 8'h1E},
{8'h03, 8'h03, 8'h19},
{8'h01, 8'h00, 8'h0F},
{8'h2F, 8'h2F, 8'h36},
{8'h80, 8'h7E, 8'h82},
{8'h80, 8'h7E, 8'h7F},
{8'h77, 8'h74, 8'h75},
{8'hA4, 8'hA0, 8'hA1},
{8'hF9, 8'hF9, 8'hF3},
{8'hF4, 8'hF4, 8'hF0},
{8'h90, 8'h8F, 8'h8F},
{8'h7C, 8'h7A, 8'h7D},
{8'h7D, 8'h7B, 8'h7E},
{8'h7D, 8'h7C, 8'h7B},
{8'h8A, 8'h89, 8'h85},
{8'hD1, 8'hD1, 8'hCB},
{8'hA5, 8'hA3, 8'hA4},
{8'h7A, 8'h78, 8'h7A},
{8'h82, 8'h80, 8'h81},
{8'h7D, 8'h7C, 8'h7C},
{8'h7C, 8'h7B, 8'h7B},
{8'h76, 8'h74, 8'h75},
{8'h7D, 8'h7B, 8'h7C},
{8'h81, 8'h7F, 8'h80},
{8'h7F, 8'h7D, 8'h82},
{8'h7E, 8'h7C, 8'h80},
{8'h7B, 8'h79, 8'h7C},
{8'h89, 8'h87, 8'h89},
{8'hEB, 8'hEA, 8'hE9},
{8'hFA, 8'hF9, 8'hF7},
{8'hDB, 8'hDA, 8'hD7},
{8'h84, 8'h83, 8'h7F},
{8'h81, 8'h80, 8'h7B},
{8'h79, 8'h78, 8'h75},
{8'h97, 8'h96, 8'h94},
{8'hB1, 8'hB0, 8'hAF},
{8'h82, 8'h7F, 8'h82},
{8'h7E, 8'h7C, 8'h7F},
{8'h7F, 8'h7D, 8'h81},
{8'h7F, 8'h7D, 8'h82}
};

always_comb
begin
	if (left)
    CharacterRGB = ROM_Data[Address];
	else
	 CharacterRGB = Batt_rom[Address];
end

endmodule
