module three_display (
    input logic [11:0] Address,
    output logic [23:0] CharacterRGB
);



logic [23:0] ROM_Data [4095:0] = '{
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hF3, 8'hF3, 8'hF3},
{8'hEA, 8'hEA, 8'hEA},
{8'hEA, 8'hEA, 8'hEA},
{8'hED, 8'hED, 8'hED},
{8'hEB, 8'hEB, 8'hEB},
{8'hEA, 8'hEA, 8'hEA},
{8'hED, 8'hED, 8'hED},
{8'hEB, 8'hEB, 8'hEB},
{8'hEA, 8'hEA, 8'hEA},
{8'hEC, 8'hEC, 8'hEC},
{8'hEC, 8'hEC, 8'hEC},
{8'hEA, 8'hEA, 8'hEA},
{8'hEB, 8'hEB, 8'hEB},
{8'hED, 8'hED, 8'hED},
{8'hEA, 8'hEA, 8'hEA},
{8'hEA, 8'hEA, 8'hEA},
{8'hED, 8'hED, 8'hED},
{8'hEA, 8'hEA, 8'hEA},
{8'hEA, 8'hEA, 8'hEA},
{8'hF3, 8'hF3, 8'hF3},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'h7D, 8'h7D, 8'h7D},
{8'h15, 8'h15, 8'h15},
{8'h15, 8'h15, 8'h15},
{8'h3A, 8'h3A, 8'h3A},
{8'h17, 8'h17, 8'h17},
{8'h15, 8'h15, 8'h15},
{8'h34, 8'h34, 8'h34},
{8'h20, 8'h20, 8'h20},
{8'h15, 8'h15, 8'h15},
{8'h2A, 8'h2A, 8'h2A},
{8'h2A, 8'h2A, 8'h2A},
{8'h15, 8'h15, 8'h15},
{8'h20, 8'h20, 8'h20},
{8'h34, 8'h34, 8'h34},
{8'h15, 8'h15, 8'h15},
{8'h17, 8'h17, 8'h17},
{8'h3A, 8'h3A, 8'h3A},
{8'h15, 8'h15, 8'h15},
{8'h15, 8'h15, 8'h15},
{8'h7D, 8'h7D, 8'h7D},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'h6F, 8'h6F, 8'h6F},
{8'h00, 8'h00, 8'h00},
{8'h00, 8'h00, 8'h00},
{8'h24, 8'h24, 8'h24},
{8'h00, 8'h00, 8'h00},
{8'h00, 8'h00, 8'h00},
{8'h1E, 8'h1E, 8'h1E},
{8'h07, 8'h07, 8'h07},
{8'h00, 8'h00, 8'h00},
{8'h12, 8'h12, 8'h12},
{8'h12, 8'h12, 8'h12},
{8'h00, 8'h00, 8'h00},
{8'h07, 8'h07, 8'h07},
{8'h1E, 8'h1E, 8'h1E},
{8'h00, 8'h00, 8'h00},
{8'h00, 8'h00, 8'h00},
{8'h24, 8'h24, 8'h24},
{8'h00, 8'h00, 8'h00},
{8'h00, 8'h00, 8'h00},
{8'h6F, 8'h6F, 8'h6F},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'h7B, 8'h7B, 8'h7B},
{8'h0F, 8'h0F, 8'h0F},
{8'h10, 8'h10, 8'h10},
{8'h35, 8'h35, 8'h35},
{8'h12, 8'h12, 8'h12},
{8'h10, 8'h10, 8'h10},
{8'h30, 8'h30, 8'h30},
{8'h1B, 8'h1B, 8'h1B},
{8'h10, 8'h10, 8'h10},
{8'h25, 8'h25, 8'h25},
{8'h25, 8'h25, 8'h25},
{8'h10, 8'h10, 8'h10},
{8'h1B, 8'h1B, 8'h1B},
{8'h30, 8'h30, 8'h30},
{8'h10, 8'h10, 8'h10},
{8'h12, 8'h12, 8'h12},
{8'h35, 8'h35, 8'h35},
{8'h10, 8'h10, 8'h10},
{8'h0F, 8'h0F, 8'h0F},
{8'h7B, 8'h7B, 8'h7B},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'h6B, 8'h6B, 8'h6B},
{8'h39, 8'h39, 8'h39},
{8'h3D, 8'h3D, 8'h3D},
{8'h48, 8'h48, 8'h48},
{8'h1E, 8'h1E, 8'h1E},
{8'h1E, 8'h1E, 8'h1E},
{8'h41, 8'h41, 8'h41},
{8'h20, 8'h20, 8'h20},
{8'h1E, 8'h1E, 8'h1E},
{8'h3C, 8'h3C, 8'h3C},
{8'h29, 8'h29, 8'h29},
{8'h1E, 8'h1E, 8'h1E},
{8'h32, 8'h32, 8'h32},
{8'h32, 8'h32, 8'h32},
{8'h1E, 8'h1E, 8'h1E},
{8'h29, 8'h29, 8'h29},
{8'h3C, 8'h3C, 8'h3C},
{8'h1E, 8'h1E, 8'h1E},
{8'h20, 8'h20, 8'h20},
{8'h42, 8'h42, 8'h42},
{8'h1E, 8'h1E, 8'h1E},
{8'h1E, 8'h1E, 8'h1E},
{8'h49, 8'h49, 8'h49},
{8'h3D, 8'h3D, 8'h3D},
{8'h39, 8'h39, 8'h39},
{8'h6A, 8'h6A, 8'h6A},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'h39, 8'h39, 8'h39},
{8'h00, 8'h00, 8'h00},
{8'h00, 8'h00, 8'h00},
{8'h22, 8'h22, 8'h22},
{8'h00, 8'h00, 8'h00},
{8'h00, 8'h00, 8'h00},
{8'h25, 8'h25, 8'h25},
{8'h00, 8'h00, 8'h00},
{8'h00, 8'h00, 8'h00},
{8'h1F, 8'h1F, 8'h1F},
{8'h09, 8'h09, 8'h09},
{8'h00, 8'h00, 8'h00},
{8'h14, 8'h14, 8'h14},
{8'h14, 8'h14, 8'h14},
{8'h00, 8'h00, 8'h00},
{8'h09, 8'h09, 8'h09},
{8'h1F, 8'h1F, 8'h1F},
{8'h00, 8'h00, 8'h00},
{8'h00, 8'h00, 8'h00},
{8'h25, 8'h25, 8'h25},
{8'h00, 8'h00, 8'h00},
{8'h00, 8'h00, 8'h00},
{8'h23, 8'h23, 8'h23},
{8'h00, 8'h00, 8'h00},
{8'h00, 8'h00, 8'h00},
{8'h39, 8'h39, 8'h39},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'h44, 8'h44, 8'h44},
{8'h05, 8'h05, 8'h05},
{8'h09, 8'h09, 8'h09},
{8'h2B, 8'h2B, 8'h2B},
{8'h05, 8'h05, 8'h05},
{8'h05, 8'h05, 8'h05},
{8'h29, 8'h29, 8'h29},
{8'h00, 8'h00, 8'h00},
{8'h00, 8'h00, 8'h00},
{8'h1E, 8'h1E, 8'h1E},
{8'h08, 8'h08, 8'h08},
{8'h00, 8'h00, 8'h00},
{8'h13, 8'h13, 8'h13},
{8'h13, 8'h13, 8'h13},
{8'h00, 8'h00, 8'h00},
{8'h08, 8'h08, 8'h08},
{8'h1E, 8'h1E, 8'h1E},
{8'h00, 8'h00, 8'h00},
{8'h00, 8'h00, 8'h00},
{8'h29, 8'h29, 8'h29},
{8'h05, 8'h05, 8'h05},
{8'h05, 8'h05, 8'h05},
{8'h2B, 8'h2B, 8'h2B},
{8'h09, 8'h09, 8'h09},
{8'h05, 8'h05, 8'h05},
{8'h44, 8'h44, 8'h44},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hF5, 8'hF5, 8'hF5},
{8'h78, 8'h78, 8'h78},
{8'h69, 8'h69, 8'h69},
{8'h73, 8'h73, 8'h73},
{8'h49, 8'h49, 8'h49},
{8'h25, 8'h25, 8'h25},
{8'h29, 8'h29, 8'h29},
{8'h46, 8'h46, 8'h46},
{8'h25, 8'h25, 8'h25},
{8'h25, 8'h25, 8'h25},
{8'h7B, 8'h7B, 8'h7B},
{8'hBB, 8'hBB, 8'hBB},
{8'hBA, 8'hBA, 8'hBA},
{8'hC3, 8'hC3, 8'hC3},
{8'hBE, 8'hBE, 8'hBE},
{8'hBA, 8'hBA, 8'hBA},
{8'hC0, 8'hC0, 8'hC0},
{8'hC0, 8'hC0, 8'hC0},
{8'hBA, 8'hBA, 8'hBA},
{8'hBE, 8'hBE, 8'hBE},
{8'hC3, 8'hC3, 8'hC3},
{8'hBA, 8'hBA, 8'hBA},
{8'hBB, 8'hBB, 8'hBB},
{8'h7C, 8'h7C, 8'h7C},
{8'h25, 8'h25, 8'h25},
{8'h25, 8'h25, 8'h25},
{8'h47, 8'h47, 8'h47},
{8'h29, 8'h29, 8'h29},
{8'h25, 8'h25, 8'h25},
{8'h49, 8'h49, 8'h49},
{8'h73, 8'h73, 8'h73},
{8'h69, 8'h69, 8'h69},
{8'h78, 8'h78, 8'h78},
{8'hF4, 8'hF4, 8'hF4},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hED, 8'hED, 8'hED},
{8'h10, 8'h10, 8'h10},
{8'h00, 8'h00, 8'h00},
{8'h05, 8'h05, 8'h05},
{8'h1C, 8'h1C, 8'h1C},
{8'h00, 8'h00, 8'h00},
{8'h02, 8'h02, 8'h02},
{8'h24, 8'h24, 8'h24},
{8'h00, 8'h00, 8'h00},
{8'h00, 8'h00, 8'h00},
{8'h83, 8'h83, 8'h83},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'h83, 8'h83, 8'h83},
{8'h00, 8'h00, 8'h00},
{8'h00, 8'h00, 8'h00},
{8'h25, 8'h25, 8'h25},
{8'h02, 8'h02, 8'h02},
{8'h00, 8'h00, 8'h00},
{8'h1C, 8'h1C, 8'h1C},
{8'h05, 8'h05, 8'h05},
{8'h00, 8'h00, 8'h00},
{8'h0F, 8'h0F, 8'h0F},
{8'hEC, 8'hEC, 8'hEC},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hEE, 8'hEE, 8'hEE},
{8'h18, 8'h18, 8'h18},
{8'h00, 8'h00, 8'h00},
{8'h0E, 8'h0E, 8'h0E},
{8'h1E, 8'h1E, 8'h1E},
{8'h00, 8'h00, 8'h00},
{8'h03, 8'h03, 8'h03},
{8'h20, 8'h20, 8'h20},
{8'h00, 8'h00, 8'h00},
{8'h00, 8'h00, 8'h00},
{8'h7C, 8'h7C, 8'h7C},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'h7C, 8'h7C, 8'h7C},
{8'h00, 8'h00, 8'h00},
{8'h00, 8'h00, 8'h00},
{8'h21, 8'h21, 8'h21},
{8'h03, 8'h03, 8'h03},
{8'h00, 8'h00, 8'h00},
{8'h1E, 8'h1E, 8'h1E},
{8'h0E, 8'h0E, 8'h0E},
{8'h00, 8'h00, 8'h00},
{8'h17, 8'h17, 8'h17},
{8'hED, 8'hED, 8'hED},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hF1, 8'hF1, 8'hF1},
{8'h3D, 8'h3D, 8'h3D},
{8'h27, 8'h27, 8'h27},
{8'h35, 8'h35, 8'h35},
{8'h43, 8'h43, 8'h43},
{8'h28, 8'h28, 8'h28},
{8'h2A, 8'h2A, 8'h2A},
{8'h7C, 8'h7C, 8'h7C},
{8'h87, 8'h87, 8'h87},
{8'h86, 8'h86, 8'h86},
{8'hC3, 8'hC3, 8'hC3},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hC3, 8'hC3, 8'hC3},
{8'h86, 8'h86, 8'h86},
{8'h87, 8'h87, 8'h87},
{8'h7D, 8'h7D, 8'h7D},
{8'h2A, 8'h2A, 8'h2A},
{8'h28, 8'h28, 8'h28},
{8'h43, 8'h43, 8'h43},
{8'h35, 8'h35, 8'h35},
{8'h27, 8'h27, 8'h27},
{8'h3D, 8'h3D, 8'h3D},
{8'hF0, 8'hF0, 8'hF0},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hEE, 8'hEE, 8'hEE},
{8'h1A, 8'h1A, 8'h1A},
{8'h01, 8'h01, 8'h01},
{8'h10, 8'h10, 8'h10},
{8'h20, 8'h20, 8'h20},
{8'h01, 8'h01, 8'h01},
{8'h01, 8'h01, 8'h01},
{8'hB9, 8'hB9, 8'hB9},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hB9, 8'hB9, 8'hB9},
{8'h01, 8'h01, 8'h01},
{8'h01, 8'h01, 8'h01},
{8'h20, 8'h20, 8'h20},
{8'h10, 8'h10, 8'h10},
{8'h01, 8'h01, 8'h01},
{8'h1A, 8'h1A, 8'h1A},
{8'hED, 8'hED, 8'hED},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hEE, 8'hEE, 8'hEE},
{8'h16, 8'h16, 8'h16},
{8'h00, 8'h00, 8'h00},
{8'h0C, 8'h0C, 8'h0C},
{8'h1C, 8'h1C, 8'h1C},
{8'h00, 8'h00, 8'h00},
{8'h00, 8'h00, 8'h00},
{8'hB2, 8'hB2, 8'hB2},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hB0, 8'hB0, 8'hB0},
{8'h00, 8'h00, 8'h00},
{8'h00, 8'h00, 8'h00},
{8'h17, 8'h17, 8'h17},
{8'h06, 8'h06, 8'h06},
{8'h00, 8'h00, 8'h00},
{8'h10, 8'h10, 8'h10},
{8'hEC, 8'hEC, 8'hEC},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hF0, 8'hF0, 8'hF0},
{8'h39, 8'h39, 8'h39},
{8'h23, 8'h23, 8'h23},
{8'h30, 8'h30, 8'h30},
{8'h3E, 8'h3E, 8'h3E},
{8'h23, 8'h23, 8'h23},
{8'h23, 8'h23, 8'h23},
{8'hBD, 8'hBD, 8'hBD},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hCC, 8'hCC, 8'hCC},
{8'h53, 8'h53, 8'h53},
{8'h53, 8'h53, 8'h53},
{8'h68, 8'h68, 8'h68},
{8'h5D, 8'h5D, 8'h5D},
{8'h53, 8'h53, 8'h53},
{8'h63, 8'h63, 8'h63},
{8'hF3, 8'hF3, 8'hF3},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hEF, 8'hEF, 8'hEF},
{8'h22, 8'h22, 8'h22},
{8'h0A, 8'h0A, 8'h0A},
{8'h18, 8'h18, 8'h18},
{8'h28, 8'h28, 8'h28},
{8'h0A, 8'h0A, 8'h0A},
{8'h0A, 8'h0A, 8'h0A},
{8'hB6, 8'hB6, 8'hB6},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hEE, 8'hEE, 8'hEE},
{8'h16, 8'h16, 8'h16},
{8'h00, 8'h00, 8'h00},
{8'h0B, 8'h0B, 8'h0B},
{8'h1C, 8'h1C, 8'h1C},
{8'h00, 8'h00, 8'h00},
{8'h00, 8'h00, 8'h00},
{8'hB3, 8'hB3, 8'hB3},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hEF, 8'hEF, 8'hEF},
{8'h30, 8'h30, 8'h30},
{8'h19, 8'h19, 8'h19},
{8'h27, 8'h27, 8'h27},
{8'h36, 8'h36, 8'h36},
{8'h19, 8'h19, 8'h19},
{8'h1A, 8'h1A, 8'h1A},
{8'hB3, 8'hB3, 8'hB3},
{8'hF2, 8'hF2, 8'hF2},
{8'hF1, 8'hF1, 8'hF1},
{8'hF8, 8'hF8, 8'hF8},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hEF, 8'hEF, 8'hEF},
{8'h2D, 8'h2D, 8'h2D},
{8'h16, 8'h16, 8'h16},
{8'h24, 8'h24, 8'h24},
{8'h33, 8'h33, 8'h33},
{8'h16, 8'h16, 8'h16},
{8'h1A, 8'h1A, 8'h1A},
{8'h3D, 8'h3D, 8'h3D},
{8'h1D, 8'h1D, 8'h1D},
{8'h1D, 8'h1D, 8'h1D},
{8'h8F, 8'h8F, 8'h8F},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hEE, 8'hEE, 8'hEE},
{8'h15, 8'h15, 8'h15},
{8'h00, 8'h00, 8'h00},
{8'h0B, 8'h0B, 8'h0B},
{8'h1B, 8'h1B, 8'h1B},
{8'h00, 8'h00, 8'h00},
{8'h00, 8'h00, 8'h00},
{8'h22, 8'h22, 8'h22},
{8'h00, 8'h00, 8'h00},
{8'h00, 8'h00, 8'h00},
{8'h7E, 8'h7E, 8'h7E},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hEE, 8'hEE, 8'hEE},
{8'h20, 8'h20, 8'h20},
{8'h08, 8'h08, 8'h08},
{8'h16, 8'h16, 8'h16},
{8'h2A, 8'h2A, 8'h2A},
{8'h0D, 8'h0D, 8'h0D},
{8'h11, 8'h11, 8'h11},
{8'h31, 8'h31, 8'h31},
{8'h0D, 8'h0D, 8'h0D},
{8'h0C, 8'h0C, 8'h0C},
{8'h89, 8'h89, 8'h89},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFC, 8'hFC, 8'hFC},
{8'hDD, 8'hDD, 8'hDD},
{8'hD9, 8'hD9, 8'hD9},
{8'hDC, 8'hDC, 8'hDC},
{8'h53, 8'h53, 8'h53},
{8'h20, 8'h20, 8'h20},
{8'h25, 8'h25, 8'h25},
{8'h42, 8'h42, 8'h42},
{8'h20, 8'h20, 8'h20},
{8'h20, 8'h20, 8'h20},
{8'h51, 8'h51, 8'h51},
{8'h48, 8'h48, 8'h48},
{8'h46, 8'h46, 8'h46},
{8'h5F, 8'h5F, 8'h5F},
{8'h4F, 8'h4F, 8'h4F},
{8'h46, 8'h46, 8'h46},
{8'h57, 8'h57, 8'h57},
{8'h57, 8'h57, 8'h57},
{8'h46, 8'h46, 8'h46},
{8'h4F, 8'h4F, 8'h4F},
{8'h5F, 8'h5F, 8'h5F},
{8'h46, 8'h46, 8'h46},
{8'h46, 8'h46, 8'h46},
{8'hBF, 8'hBF, 8'hBF},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'h3D, 8'h3D, 8'h3D},
{8'h00, 8'h00, 8'h00},
{8'h01, 8'h01, 8'h01},
{8'h23, 8'h23, 8'h23},
{8'h00, 8'h00, 8'h00},
{8'h00, 8'h00, 8'h00},
{8'h24, 8'h24, 8'h24},
{8'h00, 8'h00, 8'h00},
{8'h00, 8'h00, 8'h00},
{8'h1B, 8'h1B, 8'h1B},
{8'h04, 8'h04, 8'h04},
{8'h00, 8'h00, 8'h00},
{8'h0F, 8'h0F, 8'h0F},
{8'h0F, 8'h0F, 8'h0F},
{8'h00, 8'h00, 8'h00},
{8'h04, 8'h04, 8'h04},
{8'h1B, 8'h1B, 8'h1B},
{8'h00, 8'h00, 8'h00},
{8'h00, 8'h00, 8'h00},
{8'hA3, 8'hA3, 8'hA3},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'h42, 8'h42, 8'h42},
{8'h03, 8'h03, 8'h03},
{8'h07, 8'h07, 8'h07},
{8'h29, 8'h29, 8'h29},
{8'h03, 8'h03, 8'h03},
{8'h03, 8'h03, 8'h03},
{8'h2B, 8'h2B, 8'h2B},
{8'h05, 8'h05, 8'h05},
{8'h03, 8'h03, 8'h03},
{8'h25, 8'h25, 8'h25},
{8'h0F, 8'h0F, 8'h0F},
{8'h03, 8'h03, 8'h03},
{8'h1A, 8'h1A, 8'h1A},
{8'h1A, 8'h1A, 8'h1A},
{8'h03, 8'h03, 8'h03},
{8'h0F, 8'h0F, 8'h0F},
{8'h25, 8'h25, 8'h25},
{8'h03, 8'h03, 8'h03},
{8'h03, 8'h03, 8'h03},
{8'hA7, 8'hA7, 8'hA7},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'h5D, 8'h5D, 8'h5D},
{8'h26, 8'h26, 8'h26},
{8'h2B, 8'h2B, 8'h2B},
{8'h48, 8'h48, 8'h48},
{8'h27, 8'h27, 8'h27},
{8'h27, 8'h27, 8'h27},
{8'h49, 8'h49, 8'h49},
{8'h2A, 8'h2A, 8'h2A},
{8'h27, 8'h27, 8'h27},
{8'h44, 8'h44, 8'h44},
{8'h32, 8'h32, 8'h32},
{8'h27, 8'h27, 8'h27},
{8'h3B, 8'h3B, 8'h3B},
{8'h3B, 8'h3B, 8'h3B},
{8'h27, 8'h27, 8'h27},
{8'h32, 8'h32, 8'h32},
{8'h44, 8'h44, 8'h44},
{8'h27, 8'h27, 8'h27},
{8'h26, 8'h26, 8'h26},
{8'hB4, 8'hB4, 8'hB4},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'h3E, 8'h3E, 8'h3E},
{8'h00, 8'h00, 8'h00},
{8'h02, 8'h02, 8'h02},
{8'h25, 8'h25, 8'h25},
{8'h00, 8'h00, 8'h00},
{8'h00, 8'h00, 8'h00},
{8'h27, 8'h27, 8'h27},
{8'h00, 8'h00, 8'h00},
{8'h00, 8'h00, 8'h00},
{8'h21, 8'h21, 8'h21},
{8'h0A, 8'h0A, 8'h0A},
{8'h00, 8'h00, 8'h00},
{8'h16, 8'h16, 8'h16},
{8'h16, 8'h16, 8'h16},
{8'h00, 8'h00, 8'h00},
{8'h0A, 8'h0A, 8'h0A},
{8'h21, 8'h21, 8'h21},
{8'h00, 8'h00, 8'h00},
{8'h00, 8'h00, 8'h00},
{8'hA5, 8'hA5, 8'hA5},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'h3F, 8'h3F, 8'h3F},
{8'h00, 8'h00, 8'h00},
{8'h02, 8'h02, 8'h02},
{8'h25, 8'h25, 8'h25},
{8'h00, 8'h00, 8'h00},
{8'h00, 8'h00, 8'h00},
{8'h24, 8'h24, 8'h24},
{8'h00, 8'h00, 8'h00},
{8'h00, 8'h00, 8'h00},
{8'h19, 8'h19, 8'h19},
{8'h02, 8'h02, 8'h02},
{8'h00, 8'h00, 8'h00},
{8'h0D, 8'h0D, 8'h0D},
{8'h0D, 8'h0D, 8'h0D},
{8'h00, 8'h00, 8'h00},
{8'h02, 8'h02, 8'h02},
{8'h19, 8'h19, 8'h19},
{8'h00, 8'h00, 8'h00},
{8'h00, 8'h00, 8'h00},
{8'hA2, 8'hA2, 8'hA2},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hF9, 8'hF9, 8'hF9},
{8'hB5, 8'hB5, 8'hB5},
{8'hAD, 8'hAD, 8'hAD},
{8'hB2, 8'hB2, 8'hB2},
{8'h52, 8'h52, 8'h52},
{8'h27, 8'h27, 8'h27},
{8'h2B, 8'h2B, 8'h2B},
{8'h48, 8'h48, 8'h48},
{8'h27, 8'h27, 8'h27},
{8'h27, 8'h27, 8'h27},
{8'h65, 8'h65, 8'h65},
{8'h7A, 8'h7A, 8'h7A},
{8'h78, 8'h78, 8'h78},
{8'h8A, 8'h8A, 8'h8A},
{8'h7F, 8'h7F, 8'h7F},
{8'h78, 8'h78, 8'h78},
{8'h84, 8'h84, 8'h84},
{8'h84, 8'h84, 8'h84},
{8'h78, 8'h78, 8'h78},
{8'h7E, 8'h7E, 8'h7E},
{8'h8A, 8'h8A, 8'h8A},
{8'h78, 8'h78, 8'h78},
{8'h78, 8'h78, 8'h78},
{8'hD0, 8'hD0, 8'hD0},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hED, 8'hED, 8'hED},
{8'h12, 8'h12, 8'h12},
{8'h00, 8'h00, 8'h00},
{8'h08, 8'h08, 8'h08},
{8'h21, 8'h21, 8'h21},
{8'h03, 8'h03, 8'h03},
{8'h07, 8'h07, 8'h07},
{8'h29, 8'h29, 8'h29},
{8'h03, 8'h03, 8'h03},
{8'h03, 8'h03, 8'h03},
{8'h86, 8'h86, 8'h86},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hEE, 8'hEE, 8'hEE},
{8'h16, 8'h16, 8'h16},
{8'h00, 8'h00, 8'h00},
{8'h0C, 8'h0C, 8'h0C},
{8'h1C, 8'h1C, 8'h1C},
{8'h00, 8'h00, 8'h00},
{8'h01, 8'h01, 8'h01},
{8'h20, 8'h20, 8'h20},
{8'h00, 8'h00, 8'h00},
{8'h00, 8'h00, 8'h00},
{8'h7D, 8'h7D, 8'h7D},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hF0, 8'hF0, 8'hF0},
{8'h36, 8'h36, 8'h36},
{8'h20, 8'h20, 8'h20},
{8'h2E, 8'h2E, 8'h2E},
{8'h3C, 8'h3C, 8'h3C},
{8'h20, 8'h20, 8'h20},
{8'h23, 8'h23, 8'h23},
{8'h56, 8'h56, 8'h56},
{8'h46, 8'h46, 8'h46},
{8'h45, 8'h45, 8'h45},
{8'hA3, 8'hA3, 8'hA3},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hEF, 8'hEF, 8'hEF},
{8'h24, 8'h24, 8'h24},
{8'h0D, 8'h0D, 8'h0D},
{8'h1B, 8'h1B, 8'h1B},
{8'h2A, 8'h2A, 8'h2A},
{8'h0D, 8'h0D, 8'h0D},
{8'h0D, 8'h0D, 8'h0D},
{8'hB9, 8'hB9, 8'hB9},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hEE, 8'hEE, 8'hEE},
{8'h16, 8'h16, 8'h16},
{8'h00, 8'h00, 8'h00},
{8'h0B, 8'h0B, 8'h0B},
{8'h1C, 8'h1C, 8'h1C},
{8'h00, 8'h00, 8'h00},
{8'h00, 8'h00, 8'h00},
{8'hB2, 8'hB2, 8'hB2},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hEF, 8'hEF, 8'hEF},
{8'h2D, 8'h2D, 8'h2D},
{8'h16, 8'h16, 8'h16},
{8'h24, 8'h24, 8'h24},
{8'h33, 8'h33, 8'h33},
{8'h16, 8'h16, 8'h16},
{8'h16, 8'h16, 8'h16},
{8'hBA, 8'hBA, 8'hBA},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hF0, 8'hF0, 8'hF0},
{8'h30, 8'h30, 8'h30},
{8'h19, 8'h19, 8'h19},
{8'h27, 8'h27, 8'h27},
{8'h35, 8'h35, 8'h35},
{8'h19, 8'h19, 8'h19},
{8'h19, 8'h19, 8'h19},
{8'hBA, 8'hBA, 8'hBA},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hEE, 8'hEE, 8'hEE},
{8'h16, 8'h16, 8'h16},
{8'h00, 8'h00, 8'h00},
{8'h0B, 8'h0B, 8'h0B},
{8'h1C, 8'h1C, 8'h1C},
{8'h00, 8'h00, 8'h00},
{8'h00, 8'h00, 8'h00},
{8'hB2, 8'hB2, 8'hB2},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hEF, 8'hEF, 8'hEF},
{8'h22, 8'h22, 8'h22},
{8'h0A, 8'h0A, 8'h0A},
{8'h19, 8'h19, 8'h19},
{8'h28, 8'h28, 8'h28},
{8'h0A, 8'h0A, 8'h0A},
{8'h0A, 8'h0A, 8'h0A},
{8'hB6, 8'hB6, 8'hB6},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hF0, 8'hF0, 8'hF0},
{8'h39, 8'h39, 8'h39},
{8'h23, 8'h23, 8'h23},
{8'h30, 8'h30, 8'h30},
{8'h3E, 8'h3E, 8'h3E},
{8'h23, 8'h23, 8'h23},
{8'h23, 8'h23, 8'h23},
{8'hBD, 8'hBD, 8'hBD},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hCC, 8'hCC, 8'hCC},
{8'h53, 8'h53, 8'h53},
{8'h53, 8'h53, 8'h53},
{8'h68, 8'h68, 8'h68},
{8'h5D, 8'h5D, 8'h5D},
{8'h53, 8'h53, 8'h53},
{8'h63, 8'h63, 8'h63},
{8'hF3, 8'hF3, 8'hF3},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hEE, 8'hEE, 8'hEE},
{8'h16, 8'h16, 8'h16},
{8'h00, 8'h00, 8'h00},
{8'h0C, 8'h0C, 8'h0C},
{8'h1C, 8'h1C, 8'h1C},
{8'h00, 8'h00, 8'h00},
{8'h00, 8'h00, 8'h00},
{8'hB2, 8'hB2, 8'hB2},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hB0, 8'hB0, 8'hB0},
{8'h00, 8'h00, 8'h00},
{8'h00, 8'h00, 8'h00},
{8'h17, 8'h17, 8'h17},
{8'h06, 8'h06, 8'h06},
{8'h00, 8'h00, 8'h00},
{8'h10, 8'h10, 8'h10},
{8'hEC, 8'hEC, 8'hEC},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hEE, 8'hEE, 8'hEE},
{8'h1A, 8'h1A, 8'h1A},
{8'h01, 8'h01, 8'h01},
{8'h10, 8'h10, 8'h10},
{8'h21, 8'h21, 8'h21},
{8'h01, 8'h01, 8'h01},
{8'h01, 8'h01, 8'h01},
{8'hB9, 8'hB9, 8'hB9},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hB9, 8'hB9, 8'hB9},
{8'h01, 8'h01, 8'h01},
{8'h01, 8'h01, 8'h01},
{8'h20, 8'h20, 8'h20},
{8'h11, 8'h11, 8'h11},
{8'h01, 8'h01, 8'h01},
{8'h1A, 8'h1A, 8'h1A},
{8'hED, 8'hED, 8'hED},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hF0, 8'hF0, 8'hF0},
{8'h3E, 8'h3E, 8'h3E},
{8'h28, 8'h28, 8'h28},
{8'h35, 8'h35, 8'h35},
{8'h43, 8'h43, 8'h43},
{8'h28, 8'h28, 8'h28},
{8'h2A, 8'h2A, 8'h2A},
{8'h7D, 8'h7D, 8'h7D},
{8'h87, 8'h87, 8'h87},
{8'h86, 8'h86, 8'h86},
{8'hC3, 8'hC3, 8'hC3},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hC3, 8'hC3, 8'hC3},
{8'h86, 8'h86, 8'h86},
{8'h87, 8'h87, 8'h87},
{8'h7D, 8'h7D, 8'h7D},
{8'h2A, 8'h2A, 8'h2A},
{8'h28, 8'h28, 8'h28},
{8'h43, 8'h43, 8'h43},
{8'h35, 8'h35, 8'h35},
{8'h28, 8'h28, 8'h28},
{8'h3D, 8'h3D, 8'h3D},
{8'hF0, 8'hF0, 8'hF0},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hEE, 8'hEE, 8'hEE},
{8'h18, 8'h18, 8'h18},
{8'h00, 8'h00, 8'h00},
{8'h0E, 8'h0E, 8'h0E},
{8'h1E, 8'h1E, 8'h1E},
{8'h00, 8'h00, 8'h00},
{8'h03, 8'h03, 8'h03},
{8'h20, 8'h20, 8'h20},
{8'h00, 8'h00, 8'h00},
{8'h00, 8'h00, 8'h00},
{8'h7C, 8'h7C, 8'h7C},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'h7C, 8'h7C, 8'h7C},
{8'h00, 8'h00, 8'h00},
{8'h00, 8'h00, 8'h00},
{8'h21, 8'h21, 8'h21},
{8'h03, 8'h03, 8'h03},
{8'h00, 8'h00, 8'h00},
{8'h1E, 8'h1E, 8'h1E},
{8'h0E, 8'h0E, 8'h0E},
{8'h00, 8'h00, 8'h00},
{8'h17, 8'h17, 8'h17},
{8'hED, 8'hED, 8'hED},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hED, 8'hED, 8'hED},
{8'h10, 8'h10, 8'h10},
{8'h00, 8'h00, 8'h00},
{8'h05, 8'h05, 8'h05},
{8'h1C, 8'h1C, 8'h1C},
{8'h00, 8'h00, 8'h00},
{8'h02, 8'h02, 8'h02},
{8'h24, 8'h24, 8'h24},
{8'h00, 8'h00, 8'h00},
{8'h00, 8'h00, 8'h00},
{8'h83, 8'h83, 8'h83},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'h83, 8'h83, 8'h83},
{8'h00, 8'h00, 8'h00},
{8'h00, 8'h00, 8'h00},
{8'h25, 8'h25, 8'h25},
{8'h02, 8'h02, 8'h02},
{8'h00, 8'h00, 8'h00},
{8'h1C, 8'h1C, 8'h1C},
{8'h05, 8'h05, 8'h05},
{8'h00, 8'h00, 8'h00},
{8'h0F, 8'h0F, 8'h0F},
{8'hEC, 8'hEC, 8'hEC},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hF5, 8'hF5, 8'hF5},
{8'h79, 8'h79, 8'h79},
{8'h69, 8'h69, 8'h69},
{8'h73, 8'h73, 8'h73},
{8'h49, 8'h49, 8'h49},
{8'h25, 8'h25, 8'h25},
{8'h29, 8'h29, 8'h29},
{8'h46, 8'h46, 8'h46},
{8'h25, 8'h25, 8'h25},
{8'h25, 8'h25, 8'h25},
{8'h7B, 8'h7B, 8'h7B},
{8'hBB, 8'hBB, 8'hBB},
{8'hBA, 8'hBA, 8'hBA},
{8'hC4, 8'hC4, 8'hC4},
{8'hBE, 8'hBE, 8'hBE},
{8'hBA, 8'hBA, 8'hBA},
{8'hC1, 8'hC1, 8'hC1},
{8'hC1, 8'hC1, 8'hC1},
{8'hBA, 8'hBA, 8'hBA},
{8'hBE, 8'hBE, 8'hBE},
{8'hC4, 8'hC4, 8'hC4},
{8'hBA, 8'hBA, 8'hBA},
{8'hBB, 8'hBB, 8'hBB},
{8'h7C, 8'h7C, 8'h7C},
{8'h25, 8'h25, 8'h25},
{8'h25, 8'h25, 8'h25},
{8'h47, 8'h47, 8'h47},
{8'h29, 8'h29, 8'h29},
{8'h25, 8'h25, 8'h25},
{8'h49, 8'h49, 8'h49},
{8'h72, 8'h72, 8'h72},
{8'h69, 8'h69, 8'h69},
{8'h78, 8'h78, 8'h78},
{8'hF5, 8'hF5, 8'hF5},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'h44, 8'h44, 8'h44},
{8'h05, 8'h05, 8'h05},
{8'h09, 8'h09, 8'h09},
{8'h2B, 8'h2B, 8'h2B},
{8'h05, 8'h05, 8'h05},
{8'h05, 8'h05, 8'h05},
{8'h29, 8'h29, 8'h29},
{8'h00, 8'h00, 8'h00},
{8'h00, 8'h00, 8'h00},
{8'h1E, 8'h1E, 8'h1E},
{8'h08, 8'h08, 8'h08},
{8'h00, 8'h00, 8'h00},
{8'h13, 8'h13, 8'h13},
{8'h13, 8'h13, 8'h13},
{8'h00, 8'h00, 8'h00},
{8'h08, 8'h08, 8'h08},
{8'h1E, 8'h1E, 8'h1E},
{8'h00, 8'h00, 8'h00},
{8'h00, 8'h00, 8'h00},
{8'h29, 8'h29, 8'h29},
{8'h05, 8'h05, 8'h05},
{8'h05, 8'h05, 8'h05},
{8'h2C, 8'h2C, 8'h2C},
{8'h09, 8'h09, 8'h09},
{8'h05, 8'h05, 8'h05},
{8'h44, 8'h44, 8'h44},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'h39, 8'h39, 8'h39},
{8'h00, 8'h00, 8'h00},
{8'h00, 8'h00, 8'h00},
{8'h22, 8'h22, 8'h22},
{8'h00, 8'h00, 8'h00},
{8'h00, 8'h00, 8'h00},
{8'h25, 8'h25, 8'h25},
{8'h00, 8'h00, 8'h00},
{8'h00, 8'h00, 8'h00},
{8'h1F, 8'h1F, 8'h1F},
{8'h09, 8'h09, 8'h09},
{8'h00, 8'h00, 8'h00},
{8'h14, 8'h14, 8'h14},
{8'h14, 8'h14, 8'h14},
{8'h00, 8'h00, 8'h00},
{8'h09, 8'h09, 8'h09},
{8'h1F, 8'h1F, 8'h1F},
{8'h00, 8'h00, 8'h00},
{8'h00, 8'h00, 8'h00},
{8'h25, 8'h25, 8'h25},
{8'h00, 8'h00, 8'h00},
{8'h00, 8'h00, 8'h00},
{8'h23, 8'h23, 8'h23},
{8'h00, 8'h00, 8'h00},
{8'h00, 8'h00, 8'h00},
{8'h39, 8'h39, 8'h39},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'h6B, 8'h6B, 8'h6B},
{8'h39, 8'h39, 8'h39},
{8'h3D, 8'h3D, 8'h3D},
{8'h48, 8'h48, 8'h48},
{8'h1D, 8'h1D, 8'h1D},
{8'h1E, 8'h1E, 8'h1E},
{8'h41, 8'h41, 8'h41},
{8'h20, 8'h20, 8'h20},
{8'h1D, 8'h1D, 8'h1D},
{8'h3C, 8'h3C, 8'h3C},
{8'h28, 8'h28, 8'h28},
{8'h1D, 8'h1D, 8'h1D},
{8'h32, 8'h32, 8'h32},
{8'h32, 8'h32, 8'h32},
{8'h1D, 8'h1D, 8'h1D},
{8'h28, 8'h28, 8'h28},
{8'h3C, 8'h3C, 8'h3C},
{8'h1D, 8'h1D, 8'h1D},
{8'h20, 8'h20, 8'h20},
{8'h41, 8'h41, 8'h41},
{8'h1E, 8'h1E, 8'h1E},
{8'h1D, 8'h1D, 8'h1D},
{8'h48, 8'h48, 8'h48},
{8'h3D, 8'h3D, 8'h3D},
{8'h39, 8'h39, 8'h39},
{8'h6B, 8'h6B, 8'h6B},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'h7B, 8'h7B, 8'h7B},
{8'h0F, 8'h0F, 8'h0F},
{8'h10, 8'h10, 8'h10},
{8'h35, 8'h35, 8'h35},
{8'h12, 8'h12, 8'h12},
{8'h10, 8'h10, 8'h10},
{8'h30, 8'h30, 8'h30},
{8'h1B, 8'h1B, 8'h1B},
{8'h10, 8'h10, 8'h10},
{8'h25, 8'h25, 8'h25},
{8'h25, 8'h25, 8'h25},
{8'h10, 8'h10, 8'h10},
{8'h1B, 8'h1B, 8'h1B},
{8'h30, 8'h30, 8'h30},
{8'h10, 8'h10, 8'h10},
{8'h12, 8'h12, 8'h12},
{8'h35, 8'h35, 8'h35},
{8'h10, 8'h10, 8'h10},
{8'h0F, 8'h0F, 8'h0F},
{8'h7B, 8'h7B, 8'h7B},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'h6F, 8'h6F, 8'h6F},
{8'h00, 8'h00, 8'h00},
{8'h00, 8'h00, 8'h00},
{8'h24, 8'h24, 8'h24},
{8'h00, 8'h00, 8'h00},
{8'h00, 8'h00, 8'h00},
{8'h1E, 8'h1E, 8'h1E},
{8'h07, 8'h07, 8'h07},
{8'h00, 8'h00, 8'h00},
{8'h12, 8'h12, 8'h12},
{8'h12, 8'h12, 8'h12},
{8'h00, 8'h00, 8'h00},
{8'h07, 8'h07, 8'h07},
{8'h1E, 8'h1E, 8'h1E},
{8'h00, 8'h00, 8'h00},
{8'h00, 8'h00, 8'h00},
{8'h24, 8'h24, 8'h24},
{8'h00, 8'h00, 8'h00},
{8'h00, 8'h00, 8'h00},
{8'h6F, 8'h6F, 8'h6F},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'h7D, 8'h7D, 8'h7D},
{8'h14, 8'h14, 8'h14},
{8'h15, 8'h15, 8'h15},
{8'h39, 8'h39, 8'h39},
{8'h16, 8'h16, 8'h16},
{8'h15, 8'h15, 8'h15},
{8'h34, 8'h34, 8'h34},
{8'h20, 8'h20, 8'h20},
{8'h15, 8'h15, 8'h15},
{8'h2A, 8'h2A, 8'h2A},
{8'h2A, 8'h2A, 8'h2A},
{8'h15, 8'h15, 8'h15},
{8'h20, 8'h20, 8'h20},
{8'h34, 8'h34, 8'h34},
{8'h15, 8'h15, 8'h15},
{8'h16, 8'h16, 8'h16},
{8'h39, 8'h39, 8'h39},
{8'h15, 8'h15, 8'h15},
{8'h14, 8'h14, 8'h14},
{8'h7D, 8'h7D, 8'h7D},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hF3, 8'hF3, 8'hF3},
{8'hEA, 8'hEA, 8'hEA},
{8'hEA, 8'hEA, 8'hEA},
{8'hED, 8'hED, 8'hED},
{8'hEA, 8'hEA, 8'hEA},
{8'hEA, 8'hEA, 8'hEA},
{8'hED, 8'hED, 8'hED},
{8'hEB, 8'hEB, 8'hEB},
{8'hEA, 8'hEA, 8'hEA},
{8'hEC, 8'hEC, 8'hEC},
{8'hEC, 8'hEC, 8'hEC},
{8'hEA, 8'hEA, 8'hEA},
{8'hEB, 8'hEB, 8'hEB},
{8'hED, 8'hED, 8'hED},
{8'hEA, 8'hEA, 8'hEA},
{8'hEA, 8'hEA, 8'hEA},
{8'hED, 8'hED, 8'hED},
{8'hEA, 8'hEA, 8'hEA},
{8'hEA, 8'hEA, 8'hEA},
{8'hF3, 8'hF3, 8'hF3},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00},
{8'hFF, 8'hD7, 8'h00}
};


    assign CharacterRGB = ROM_Data[Address];


endmodule
