// state_definitions.sv
typedef enum logic [1:0] {IDLE, PLAYING, GAME_OVER} state_t;
